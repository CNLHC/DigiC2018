module lamb100Control(
    input trigger,
    input sysRst,
    output [6:0]counter,
    output [99:0]lamb
);
carry101Counter c101C(trigger,sysRst,counter);
//====================Truthtable Variable:0====================
wire tU0U115Out;
wire tU0U117Out;
wire tU0U134Out;
wire tU0U131Out;
wire tU0U135Out;
wire tU0U114Out;
wire tU0U139Out;
wire tU0U143Out;
wire tU0U12Out;
wire tU0U110Out;
wire tU0U125Out;
wire tU0U00Out;
wire tU0U126Out;
wire tU0U140Out;
wire tU0U17Out;
wire tU0U121Out;
wire tU0U136Out;
wire tU0U113Out;
wire tU0U133Out;
wire tU0U142Out;
wire tU0U141Out;
wire tU0U13Out;
wire tU0U120Out;
wire tU0U16Out;
wire tU0U118Out;
wire tU0U137Out;
wire tU0U112Out;
wire tU0U111Out;
wire tU0U14Out;
wire tU0U10Out;
wire tU0U129Out;
wire tU0U127Out;
wire tU0U130Out;
wire tU0U132Out;
wire tU0U19Out;
wire tU0U119Out;
wire tU0U15Out;
wire tU0U138Out;
wire tU0U18Out;
wire tU0U128Out;
wire tU0U144Out;
wire tU0U116Out;
wire tU0U124Out;
wire tU0U122Out;
wire tU0U11Out;
wire tU0U123Out;
or U0U00(tU0U00Out,tU0U10Out,tU0U11Out,tU0U12Out,tU0U13Out,tU0U14Out,tU0U15Out,tU0U16Out,tU0U17Out,tU0U18Out,tU0U19Out,tU0U110Out,tU0U111Out,tU0U112Out,tU0U113Out,tU0U114Out,tU0U115Out,tU0U116Out,tU0U117Out,tU0U118Out,tU0U119Out,tU0U120Out,tU0U121Out,tU0U122Out,tU0U123Out,tU0U124Out,tU0U125Out,tU0U126Out,tU0U127Out,tU0U128Out,tU0U129Out,tU0U130Out,tU0U131Out,tU0U132Out,tU0U133Out,tU0U134Out,tU0U135Out,tU0U136Out,tU0U137Out,tU0U138Out,tU0U139Out,tU0U140Out,tU0U141Out,tU0U142Out,tU0U143Out,tU0U144Out);
and U0U10(tU0U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U0U11(tU0U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U0U12(tU0U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U0U13(tU0U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U0U14(tU0U14Out,counter[5],counter[6]);
and U0U15(tU0U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U0U16(tU0U16Out,counter[2],counter[4],counter[6]);
and U0U17(tU0U17Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U0U18(tU0U18Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U0U19(tU0U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U0U110(tU0U110Out,counter[1],~counter[2],counter[4],counter[5]);
and U0U111(tU0U111Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U0U112(tU0U112Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U0U113(tU0U113Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U0U114(tU0U114Out,counter[2],~counter[4],counter[5]);
and U0U115(tU0U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U0U116(tU0U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U0U117(tU0U117Out,~counter[1],~counter[3],counter[4],counter[5]);
and U0U118(tU0U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U0U119(tU0U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U0U120(tU0U120Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U0U121(tU0U121Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U0U122(tU0U122Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U0U123(tU0U123Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U0U124(tU0U124Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U0U125(tU0U125Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U0U126(tU0U126Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U0U127(tU0U127Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U0U128(tU0U128Out,~counter[4],~counter[5],counter[6]);
and U0U129(tU0U129Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U0U130(tU0U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U0U131(tU0U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U0U132(tU0U132Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U0U133(tU0U133Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U0U134(tU0U134Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U0U135(tU0U135Out,~counter[1],~counter[5],counter[6]);
and U0U136(tU0U136Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U0U137(tU0U137Out,counter[1],~counter[2],counter[4],counter[6]);
and U0U138(tU0U138Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U0U139(tU0U139Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U0U140(tU0U140Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U0U141(tU0U141Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U0U142(tU0U142Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U0U143(tU0U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U0U144(tU0U144Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:1====================
wire tU1U00Out;
and U1U00(tU1U00Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:2====================
wire tU2U11Out;
wire tU2U00Out;
wire tU2U10Out;
or U2U00(tU2U00Out,tU2U10Out,tU2U11Out);
and U2U10(tU2U10Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U2U11(tU2U11Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:3====================
wire tU3U15Out;
wire tU3U125Out;
wire tU3U112Out;
wire tU3U17Out;
wire tU3U114Out;
wire tU3U139Out;
wire tU3U115Out;
wire tU3U113Out;
wire tU3U00Out;
wire tU3U127Out;
wire tU3U119Out;
wire tU3U16Out;
wire tU3U11Out;
wire tU3U123Out;
wire tU3U118Out;
wire tU3U12Out;
wire tU3U110Out;
wire tU3U141Out;
wire tU3U129Out;
wire tU3U13Out;
wire tU3U135Out;
wire tU3U116Out;
wire tU3U138Out;
wire tU3U128Out;
wire tU3U132Out;
wire tU3U120Out;
wire tU3U117Out;
wire tU3U142Out;
wire tU3U140Out;
wire tU3U136Out;
wire tU3U18Out;
wire tU3U124Out;
wire tU3U122Out;
wire tU3U126Out;
wire tU3U19Out;
wire tU3U130Out;
wire tU3U137Out;
wire tU3U14Out;
wire tU3U133Out;
wire tU3U111Out;
wire tU3U134Out;
wire tU3U10Out;
wire tU3U121Out;
wire tU3U131Out;
or U3U00(tU3U00Out,tU3U10Out,tU3U11Out,tU3U12Out,tU3U13Out,tU3U14Out,tU3U15Out,tU3U16Out,tU3U17Out,tU3U18Out,tU3U19Out,tU3U110Out,tU3U111Out,tU3U112Out,tU3U113Out,tU3U114Out,tU3U115Out,tU3U116Out,tU3U117Out,tU3U118Out,tU3U119Out,tU3U120Out,tU3U121Out,tU3U122Out,tU3U123Out,tU3U124Out,tU3U125Out,tU3U126Out,tU3U127Out,tU3U128Out,tU3U129Out,tU3U130Out,tU3U131Out,tU3U132Out,tU3U133Out,tU3U134Out,tU3U135Out,tU3U136Out,tU3U137Out,tU3U138Out,tU3U139Out,tU3U140Out,tU3U141Out,tU3U142Out);
and U3U10(tU3U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U3U11(tU3U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U3U12(tU3U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U3U13(tU3U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U3U14(tU3U14Out,counter[5],counter[6]);
and U3U15(tU3U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U3U16(tU3U16Out,counter[2],counter[4],counter[6]);
and U3U17(tU3U17Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U3U18(tU3U18Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U3U19(tU3U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U3U110(tU3U110Out,counter[1],~counter[2],counter[4],counter[5]);
and U3U111(tU3U111Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U3U112(tU3U112Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U3U113(tU3U113Out,counter[2],~counter[4],counter[5]);
and U3U114(tU3U114Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U3U115(tU3U115Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U3U116(tU3U116Out,~counter[1],~counter[3],counter[4],counter[5]);
and U3U117(tU3U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U3U118(tU3U118Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U3U119(tU3U119Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U3U120(tU3U120Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U3U121(tU3U121Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U3U122(tU3U122Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U3U123(tU3U123Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U3U124(tU3U124Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U3U125(tU3U125Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U3U126(tU3U126Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U3U127(tU3U127Out,~counter[4],~counter[5],counter[6]);
and U3U128(tU3U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U3U129(tU3U129Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U3U130(tU3U130Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U3U131(tU3U131Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U3U132(tU3U132Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U3U133(tU3U133Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U3U134(tU3U134Out,~counter[1],~counter[5],counter[6]);
and U3U135(tU3U135Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U3U136(tU3U136Out,counter[1],~counter[2],counter[4],counter[6]);
and U3U137(tU3U137Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U3U138(tU3U138Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U3U139(tU3U139Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U3U140(tU3U140Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U3U141(tU3U141Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U3U142(tU3U142Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:4====================
wire tU4U11Out;
wire tU4U12Out;
wire tU4U10Out;
wire tU4U00Out;
or U4U00(tU4U00Out,tU4U10Out,tU4U11Out,tU4U12Out);
and U4U10(tU4U10Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U4U11(tU4U11Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U4U12(tU4U12Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:5====================
wire tU5U10Out;
wire tU5U12Out;
wire tU5U11Out;
wire tU5U00Out;
or U5U00(tU5U00Out,tU5U10Out,tU5U11Out,tU5U12Out);
and U5U10(tU5U10Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U5U11(tU5U11Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U5U12(tU5U12Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:6====================
wire tU6U13Out;
wire tU6U00Out;
wire tU6U11Out;
wire tU6U14Out;
wire tU6U12Out;
wire tU6U10Out;
or U6U00(tU6U00Out,tU6U10Out,tU6U11Out,tU6U12Out,tU6U13Out,tU6U14Out);
and U6U10(tU6U10Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U6U11(tU6U11Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U6U12(tU6U12Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U6U13(tU6U13Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U6U14(tU6U14Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:7====================
wire tU7U13Out;
wire tU7U10Out;
wire tU7U00Out;
wire tU7U11Out;
wire tU7U12Out;
or U7U00(tU7U00Out,tU7U10Out,tU7U11Out,tU7U12Out,tU7U13Out);
and U7U10(tU7U10Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U7U11(tU7U11Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U7U12(tU7U12Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U7U13(tU7U13Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:8====================
wire tU8U17Out;
wire tU8U114Out;
wire tU8U123Out;
wire tU8U138Out;
wire tU8U112Out;
wire tU8U118Out;
wire tU8U00Out;
wire tU8U130Out;
wire tU8U18Out;
wire tU8U110Out;
wire tU8U122Out;
wire tU8U16Out;
wire tU8U127Out;
wire tU8U125Out;
wire tU8U124Out;
wire tU8U126Out;
wire tU8U14Out;
wire tU8U12Out;
wire tU8U119Out;
wire tU8U19Out;
wire tU8U13Out;
wire tU8U129Out;
wire tU8U111Out;
wire tU8U10Out;
wire tU8U117Out;
wire tU8U116Out;
wire tU8U132Out;
wire tU8U131Out;
wire tU8U115Out;
wire tU8U120Out;
wire tU8U128Out;
wire tU8U135Out;
wire tU8U11Out;
wire tU8U113Out;
wire tU8U134Out;
wire tU8U121Out;
wire tU8U133Out;
wire tU8U15Out;
wire tU8U139Out;
wire tU8U137Out;
wire tU8U136Out;
or U8U00(tU8U00Out,tU8U10Out,tU8U11Out,tU8U12Out,tU8U13Out,tU8U14Out,tU8U15Out,tU8U16Out,tU8U17Out,tU8U18Out,tU8U19Out,tU8U110Out,tU8U111Out,tU8U112Out,tU8U113Out,tU8U114Out,tU8U115Out,tU8U116Out,tU8U117Out,tU8U118Out,tU8U119Out,tU8U120Out,tU8U121Out,tU8U122Out,tU8U123Out,tU8U124Out,tU8U125Out,tU8U126Out,tU8U127Out,tU8U128Out,tU8U129Out,tU8U130Out,tU8U131Out,tU8U132Out,tU8U133Out,tU8U134Out,tU8U135Out,tU8U136Out,tU8U137Out,tU8U138Out,tU8U139Out);
and U8U10(tU8U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U8U11(tU8U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U8U12(tU8U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U8U13(tU8U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U8U14(tU8U14Out,counter[5],counter[6]);
and U8U15(tU8U15Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U8U16(tU8U16Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U8U17(tU8U17Out,counter[2],counter[4],counter[6]);
and U8U18(tU8U18Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U8U19(tU8U19Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U8U110(tU8U110Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U8U111(tU8U111Out,counter[1],~counter[2],counter[4],counter[5]);
and U8U112(tU8U112Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U8U113(tU8U113Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U8U114(tU8U114Out,counter[2],~counter[4],counter[5]);
and U8U115(tU8U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U8U116(tU8U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U8U117(tU8U117Out,~counter[1],~counter[3],counter[4],counter[5]);
and U8U118(tU8U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U8U119(tU8U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U8U120(tU8U120Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U8U121(tU8U121Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U8U122(tU8U122Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U8U123(tU8U123Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U8U124(tU8U124Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U8U125(tU8U125Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U8U126(tU8U126Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U8U127(tU8U127Out,~counter[4],~counter[5],counter[6]);
and U8U128(tU8U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U8U129(tU8U129Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U8U130(tU8U130Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U8U131(tU8U131Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U8U132(tU8U132Out,~counter[1],~counter[5],counter[6]);
and U8U133(tU8U133Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U8U134(tU8U134Out,counter[1],~counter[2],counter[4],counter[6]);
and U8U135(tU8U135Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U8U136(tU8U136Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U8U137(tU8U137Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U8U138(tU8U138Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U8U139(tU8U139Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:9====================
wire tU9U10Out;
wire tU9U12Out;
wire tU9U11Out;
wire tU9U00Out;
wire tU9U13Out;
or U9U00(tU9U00Out,tU9U10Out,tU9U11Out,tU9U12Out,tU9U13Out);
and U9U10(tU9U10Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U9U11(tU9U11Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U9U12(tU9U12Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U9U13(tU9U13Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:10====================
wire tU10U11Out;
wire tU10U13Out;
wire tU10U14Out;
wire tU10U17Out;
wire tU10U12Out;
wire tU10U00Out;
wire tU10U10Out;
wire tU10U15Out;
wire tU10U16Out;
or U10U00(tU10U00Out,tU10U10Out,tU10U11Out,tU10U12Out,tU10U13Out,tU10U14Out,tU10U15Out,tU10U16Out,tU10U17Out);
and U10U10(tU10U10Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U10U11(tU10U11Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U10U12(tU10U12Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U10U13(tU10U13Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U10U14(tU10U14Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U10U15(tU10U15Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U10U16(tU10U16Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U10U17(tU10U17Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:11====================
wire tU11U15Out;
wire tU11U13Out;
wire tU11U12Out;
wire tU11U10Out;
wire tU11U11Out;
wire tU11U00Out;
wire tU11U14Out;
or U11U00(tU11U00Out,tU11U10Out,tU11U11Out,tU11U12Out,tU11U13Out,tU11U14Out,tU11U15Out);
and U11U10(tU11U10Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U11U11(tU11U11Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U11U12(tU11U12Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U11U13(tU11U13Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U11U14(tU11U14Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U11U15(tU11U15Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:12====================
wire tU12U10Out;
wire tU12U13Out;
wire tU12U17Out;
wire tU12U18Out;
wire tU12U19Out;
wire tU12U00Out;
wire tU12U12Out;
wire tU12U15Out;
wire tU12U14Out;
wire tU12U11Out;
wire tU12U16Out;
or U12U00(tU12U00Out,tU12U10Out,tU12U11Out,tU12U12Out,tU12U13Out,tU12U14Out,tU12U15Out,tU12U16Out,tU12U17Out,tU12U18Out,tU12U19Out);
and U12U10(tU12U10Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U12U11(tU12U11Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U12U12(tU12U12Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U12U13(tU12U13Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U12U14(tU12U14Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U12U15(tU12U15Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U12U16(tU12U16Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U12U17(tU12U17Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U12U18(tU12U18Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U12U19(tU12U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:13====================
wire tU13U10Out;
wire tU13U00Out;
wire tU13U14Out;
wire tU13U12Out;
wire tU13U16Out;
wire tU13U15Out;
wire tU13U11Out;
wire tU13U13Out;
or U13U00(tU13U00Out,tU13U10Out,tU13U11Out,tU13U12Out,tU13U13Out,tU13U14Out,tU13U15Out,tU13U16Out);
and U13U10(tU13U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U13U11(tU13U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U13U12(tU13U12Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U13U13(tU13U13Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U13U14(tU13U14Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U13U15(tU13U15Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U13U16(tU13U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:14====================
wire tU14U17Out;
wire tU14U14Out;
wire tU14U19Out;
wire tU14U15Out;
wire tU14U10Out;
wire tU14U16Out;
wire tU14U11Out;
wire tU14U13Out;
wire tU14U00Out;
wire tU14U12Out;
wire tU14U18Out;
or U14U00(tU14U00Out,tU14U10Out,tU14U11Out,tU14U12Out,tU14U13Out,tU14U14Out,tU14U15Out,tU14U16Out,tU14U17Out,tU14U18Out,tU14U19Out);
and U14U10(tU14U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U14U11(tU14U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U14U12(tU14U12Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U14U13(tU14U13Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U14U14(tU14U14Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U14U15(tU14U15Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U14U16(tU14U16Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U14U17(tU14U17Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U14U18(tU14U18Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U14U19(tU14U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:15====================
wire tU15U127Out;
wire tU15U18Out;
wire tU15U117Out;
wire tU15U134Out;
wire tU15U119Out;
wire tU15U115Out;
wire tU15U124Out;
wire tU15U126Out;
wire tU15U130Out;
wire tU15U14Out;
wire tU15U111Out;
wire tU15U128Out;
wire tU15U12Out;
wire tU15U113Out;
wire tU15U136Out;
wire tU15U133Out;
wire tU15U16Out;
wire tU15U110Out;
wire tU15U120Out;
wire tU15U129Out;
wire tU15U13Out;
wire tU15U122Out;
wire tU15U10Out;
wire tU15U11Out;
wire tU15U19Out;
wire tU15U123Out;
wire tU15U114Out;
wire tU15U125Out;
wire tU15U112Out;
wire tU15U17Out;
wire tU15U135Out;
wire tU15U118Out;
wire tU15U121Out;
wire tU15U00Out;
wire tU15U132Out;
wire tU15U131Out;
wire tU15U116Out;
wire tU15U15Out;
or U15U00(tU15U00Out,tU15U10Out,tU15U11Out,tU15U12Out,tU15U13Out,tU15U14Out,tU15U15Out,tU15U16Out,tU15U17Out,tU15U18Out,tU15U19Out,tU15U110Out,tU15U111Out,tU15U112Out,tU15U113Out,tU15U114Out,tU15U115Out,tU15U116Out,tU15U117Out,tU15U118Out,tU15U119Out,tU15U120Out,tU15U121Out,tU15U122Out,tU15U123Out,tU15U124Out,tU15U125Out,tU15U126Out,tU15U127Out,tU15U128Out,tU15U129Out,tU15U130Out,tU15U131Out,tU15U132Out,tU15U133Out,tU15U134Out,tU15U135Out,tU15U136Out);
and U15U10(tU15U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U15U11(tU15U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U15U12(tU15U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U15U13(tU15U13Out,counter[5],counter[6]);
and U15U14(tU15U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U15U15(tU15U15Out,counter[2],counter[4],counter[6]);
and U15U16(tU15U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U15U17(tU15U17Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U15U18(tU15U18Out,counter[1],~counter[2],counter[4],counter[5]);
and U15U19(tU15U19Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U15U110(tU15U110Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U15U111(tU15U111Out,counter[2],~counter[4],counter[5]);
and U15U112(tU15U112Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U15U113(tU15U113Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U15U114(tU15U114Out,~counter[1],~counter[3],counter[4],counter[5]);
and U15U115(tU15U115Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U15U116(tU15U116Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U15U117(tU15U117Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U15U118(tU15U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U15U119(tU15U119Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U15U120(tU15U120Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U15U121(tU15U121Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U15U122(tU15U122Out,~counter[4],~counter[5],counter[6]);
and U15U123(tU15U123Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U15U124(tU15U124Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U15U125(tU15U125Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U15U126(tU15U126Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U15U127(tU15U127Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U15U128(tU15U128Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U15U129(tU15U129Out,~counter[1],~counter[5],counter[6]);
and U15U130(tU15U130Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U15U131(tU15U131Out,counter[1],~counter[2],counter[4],counter[6]);
and U15U132(tU15U132Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U15U133(tU15U133Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U15U134(tU15U134Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U15U135(tU15U135Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U15U136(tU15U136Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:16====================
wire tU16U19Out;
wire tU16U16Out;
wire tU16U11Out;
wire tU16U112Out;
wire tU16U12Out;
wire tU16U113Out;
wire tU16U13Out;
wire tU16U17Out;
wire tU16U111Out;
wire tU16U15Out;
wire tU16U110Out;
wire tU16U18Out;
wire tU16U14Out;
wire tU16U00Out;
wire tU16U10Out;
or U16U00(tU16U00Out,tU16U10Out,tU16U11Out,tU16U12Out,tU16U13Out,tU16U14Out,tU16U15Out,tU16U16Out,tU16U17Out,tU16U18Out,tU16U19Out,tU16U110Out,tU16U111Out,tU16U112Out,tU16U113Out);
and U16U10(tU16U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U11(tU16U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U12(tU16U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U13(tU16U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U14(tU16U14Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U15(tU16U15Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U16U16(tU16U16Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U16U17(tU16U17Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U18(tU16U18Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U16U19(tU16U19Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U16U110(tU16U110Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U16U111(tU16U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U16U112(tU16U112Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U16U113(tU16U113Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:17====================
wire tU17U16Out;
wire tU17U17Out;
wire tU17U13Out;
wire tU17U00Out;
wire tU17U14Out;
wire tU17U11Out;
wire tU17U10Out;
wire tU17U18Out;
wire tU17U19Out;
wire tU17U110Out;
wire tU17U111Out;
wire tU17U12Out;
wire tU17U15Out;
or U17U00(tU17U00Out,tU17U10Out,tU17U11Out,tU17U12Out,tU17U13Out,tU17U14Out,tU17U15Out,tU17U16Out,tU17U17Out,tU17U18Out,tU17U19Out,tU17U110Out,tU17U111Out);
and U17U10(tU17U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U17U11(tU17U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U17U12(tU17U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U17U13(tU17U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U17U14(tU17U14Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U17U15(tU17U15Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U17U16(tU17U16Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U17U17(tU17U17Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U17U18(tU17U18Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U17U19(tU17U19Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U17U110(tU17U110Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U17U111(tU17U111Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:18====================
wire tU18U15Out;
wire tU18U111Out;
wire tU18U11Out;
wire tU18U17Out;
wire tU18U00Out;
wire tU18U13Out;
wire tU18U10Out;
wire tU18U110Out;
wire tU18U19Out;
wire tU18U14Out;
wire tU18U114Out;
wire tU18U115Out;
wire tU18U16Out;
wire tU18U112Out;
wire tU18U12Out;
wire tU18U113Out;
wire tU18U18Out;
or U18U00(tU18U00Out,tU18U10Out,tU18U11Out,tU18U12Out,tU18U13Out,tU18U14Out,tU18U15Out,tU18U16Out,tU18U17Out,tU18U18Out,tU18U19Out,tU18U110Out,tU18U111Out,tU18U112Out,tU18U113Out,tU18U114Out,tU18U115Out);
and U18U10(tU18U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U11(tU18U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U12(tU18U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U13(tU18U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U14(tU18U14Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U15(tU18U15Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U18U16(tU18U16Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U18U17(tU18U17Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U18U18(tU18U18Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U19(tU18U19Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U18U110(tU18U110Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U18U111(tU18U111Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U18U112(tU18U112Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U18U113(tU18U113Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U18U114(tU18U114Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U18U115(tU18U115Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:19====================
wire tU19U19Out;
wire tU19U13Out;
wire tU19U17Out;
wire tU19U15Out;
wire tU19U110Out;
wire tU19U14Out;
wire tU19U18Out;
wire tU19U12Out;
wire tU19U00Out;
wire tU19U16Out;
wire tU19U11Out;
wire tU19U10Out;
or U19U00(tU19U00Out,tU19U10Out,tU19U11Out,tU19U12Out,tU19U13Out,tU19U14Out,tU19U15Out,tU19U16Out,tU19U17Out,tU19U18Out,tU19U19Out,tU19U110Out);
and U19U10(tU19U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U19U11(tU19U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U19U12(tU19U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U19U13(tU19U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U19U14(tU19U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U19U15(tU19U15Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U19U16(tU19U16Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U19U17(tU19U17Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U19U18(tU19U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U19U19(tU19U19Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U19U110(tU19U110Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:20====================
wire tU20U00Out;
wire tU20U15Out;
wire tU20U13Out;
wire tU20U110Out;
wire tU20U10Out;
wire tU20U19Out;
wire tU20U112Out;
wire tU20U113Out;
wire tU20U12Out;
wire tU20U11Out;
wire tU20U14Out;
wire tU20U18Out;
wire tU20U17Out;
wire tU20U16Out;
wire tU20U111Out;
or U20U00(tU20U00Out,tU20U10Out,tU20U11Out,tU20U12Out,tU20U13Out,tU20U14Out,tU20U15Out,tU20U16Out,tU20U17Out,tU20U18Out,tU20U19Out,tU20U110Out,tU20U111Out,tU20U112Out,tU20U113Out);
and U20U10(tU20U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U11(tU20U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U12(tU20U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U13(tU20U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U20U14(tU20U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U15(tU20U15Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U16(tU20U16Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U20U17(tU20U17Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U20U18(tU20U18Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U19(tU20U19Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U20U110(tU20U110Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U20U111(tU20U111Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U20U112(tU20U112Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U20U113(tU20U113Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:21====================
wire tU21U12Out;
wire tU21U13Out;
wire tU21U17Out;
wire tU21U14Out;
wire tU21U15Out;
wire tU21U00Out;
wire tU21U10Out;
wire tU21U16Out;
wire tU21U19Out;
wire tU21U110Out;
wire tU21U11Out;
wire tU21U18Out;
or U21U00(tU21U00Out,tU21U10Out,tU21U11Out,tU21U12Out,tU21U13Out,tU21U14Out,tU21U15Out,tU21U16Out,tU21U17Out,tU21U18Out,tU21U19Out,tU21U110Out);
and U21U10(tU21U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U21U11(tU21U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U21U12(tU21U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U21U13(tU21U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U21U14(tU21U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U21U15(tU21U15Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U21U16(tU21U16Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U21U17(tU21U17Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U21U18(tU21U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U21U19(tU21U19Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U21U110(tU21U110Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:22====================
wire tU22U113Out;
wire tU22U16Out;
wire tU22U112Out;
wire tU22U12Out;
wire tU22U18Out;
wire tU22U14Out;
wire tU22U118Out;
wire tU22U110Out;
wire tU22U13Out;
wire tU22U10Out;
wire tU22U111Out;
wire tU22U116Out;
wire tU22U17Out;
wire tU22U115Out;
wire tU22U19Out;
wire tU22U00Out;
wire tU22U11Out;
wire tU22U15Out;
wire tU22U119Out;
wire tU22U117Out;
wire tU22U114Out;
or U22U00(tU22U00Out,tU22U10Out,tU22U11Out,tU22U12Out,tU22U13Out,tU22U14Out,tU22U15Out,tU22U16Out,tU22U17Out,tU22U18Out,tU22U19Out,tU22U110Out,tU22U111Out,tU22U112Out,tU22U113Out,tU22U114Out,tU22U115Out,tU22U116Out,tU22U117Out,tU22U118Out,tU22U119Out);
and U22U10(tU22U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U22U11(tU22U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U12(tU22U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U13(tU22U13Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U14(tU22U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U22U15(tU22U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U16(tU22U16Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U17(tU22U17Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U22U18(tU22U18Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U22U19(tU22U19Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U22U110(tU22U110Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U111(tU22U111Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U22U112(tU22U112Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U22U113(tU22U113Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U22U114(tU22U114Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U22U115(tU22U115Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U22U116(tU22U116Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U22U117(tU22U117Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U22U118(tU22U118Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U22U119(tU22U119Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:23====================
wire tU23U113Out;
wire tU23U11Out;
wire tU23U114Out;
wire tU23U14Out;
wire tU23U110Out;
wire tU23U13Out;
wire tU23U16Out;
wire tU23U00Out;
wire tU23U12Out;
wire tU23U10Out;
wire tU23U112Out;
wire tU23U19Out;
wire tU23U18Out;
wire tU23U15Out;
wire tU23U111Out;
wire tU23U17Out;
or U23U00(tU23U00Out,tU23U10Out,tU23U11Out,tU23U12Out,tU23U13Out,tU23U14Out,tU23U15Out,tU23U16Out,tU23U17Out,tU23U18Out,tU23U19Out,tU23U110Out,tU23U111Out,tU23U112Out,tU23U113Out,tU23U114Out);
and U23U10(tU23U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U11(tU23U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U23U12(tU23U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U23U13(tU23U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U14(tU23U14Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U23U15(tU23U15Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U16(tU23U16Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U23U17(tU23U17Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U18(tU23U18Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U19(tU23U19Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U23U110(tU23U110Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U111(tU23U111Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U23U112(tU23U112Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U23U113(tU23U113Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U23U114(tU23U114Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:24====================
wire tU24U00Out;
wire tU24U10Out;
wire tU24U112Out;
wire tU24U114Out;
wire tU24U17Out;
wire tU24U111Out;
wire tU24U120Out;
wire tU24U124Out;
wire tU24U18Out;
wire tU24U119Out;
wire tU24U14Out;
wire tU24U118Out;
wire tU24U13Out;
wire tU24U19Out;
wire tU24U113Out;
wire tU24U116Out;
wire tU24U110Out;
wire tU24U16Out;
wire tU24U123Out;
wire tU24U12Out;
wire tU24U15Out;
wire tU24U115Out;
wire tU24U121Out;
wire tU24U11Out;
wire tU24U117Out;
wire tU24U122Out;
or U24U00(tU24U00Out,tU24U10Out,tU24U11Out,tU24U12Out,tU24U13Out,tU24U14Out,tU24U15Out,tU24U16Out,tU24U17Out,tU24U18Out,tU24U19Out,tU24U110Out,tU24U111Out,tU24U112Out,tU24U113Out,tU24U114Out,tU24U115Out,tU24U116Out,tU24U117Out,tU24U118Out,tU24U119Out,tU24U120Out,tU24U121Out,tU24U122Out,tU24U123Out,tU24U124Out);
and U24U10(tU24U10Out,counter[5],counter[6]);
and U24U11(tU24U11Out,counter[2],counter[4],counter[6]);
and U24U12(tU24U12Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U24U13(tU24U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U24U14(tU24U14Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U24U15(tU24U15Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U24U16(tU24U16Out,counter[0],counter[3],counter[4],~counter[5],~counter[6]);
and U24U17(tU24U17Out,counter[2],~counter[4],counter[5]);
and U24U18(tU24U18Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U24U19(tU24U19Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U24U110(tU24U110Out,~counter[1],~counter[3],counter[4],counter[5]);
and U24U111(tU24U111Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U24U112(tU24U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U24U113(tU24U113Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U24U114(tU24U114Out,~counter[4],~counter[5],counter[6]);
and U24U115(tU24U115Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U24U116(tU24U116Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U24U117(tU24U117Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U24U118(tU24U118Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U24U119(tU24U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U24U120(tU24U120Out,~counter[1],~counter[5],counter[6]);
and U24U121(tU24U121Out,counter[1],~counter[2],counter[4],counter[6]);
and U24U122(tU24U122Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U24U123(tU24U123Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U24U124(tU24U124Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:25====================
wire tU25U111Out;
wire tU25U14Out;
wire tU25U11Out;
wire tU25U13Out;
wire tU25U19Out;
wire tU25U16Out;
wire tU25U10Out;
wire tU25U18Out;
wire tU25U00Out;
wire tU25U110Out;
wire tU25U17Out;
wire tU25U12Out;
wire tU25U15Out;
or U25U00(tU25U00Out,tU25U10Out,tU25U11Out,tU25U12Out,tU25U13Out,tU25U14Out,tU25U15Out,tU25U16Out,tU25U17Out,tU25U18Out,tU25U19Out,tU25U110Out,tU25U111Out);
and U25U10(tU25U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U11(tU25U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U25U12(tU25U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U25U13(tU25U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U14(tU25U14Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U15(tU25U15Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U16(tU25U16Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U17(tU25U17Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U25U18(tU25U18Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U19(tU25U19Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U25U110(tU25U110Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U25U111(tU25U111Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:26====================
wire tU26U112Out;
wire tU26U18Out;
wire tU26U117Out;
wire tU26U16Out;
wire tU26U115Out;
wire tU26U113Out;
wire tU26U11Out;
wire tU26U116Out;
wire tU26U12Out;
wire tU26U111Out;
wire tU26U14Out;
wire tU26U19Out;
wire tU26U114Out;
wire tU26U13Out;
wire tU26U110Out;
wire tU26U15Out;
wire tU26U00Out;
wire tU26U17Out;
wire tU26U10Out;
or U26U00(tU26U00Out,tU26U10Out,tU26U11Out,tU26U12Out,tU26U13Out,tU26U14Out,tU26U15Out,tU26U16Out,tU26U17Out,tU26U18Out,tU26U19Out,tU26U110Out,tU26U111Out,tU26U112Out,tU26U113Out,tU26U114Out,tU26U115Out,tU26U116Out,tU26U117Out);
and U26U10(tU26U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U11(tU26U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U26U12(tU26U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U26U13(tU26U13Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U26U14(tU26U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U15(tU26U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U26U16(tU26U16Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U26U17(tU26U17Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U18(tU26U18Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U19(tU26U19Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U26U110(tU26U110Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U111(tU26U111Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U26U112(tU26U112Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U113(tU26U113Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U26U114(tU26U114Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U26U115(tU26U115Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U26U116(tU26U116Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U26U117(tU26U117Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:27====================
wire tU27U115Out;
wire tU27U14Out;
wire tU27U10Out;
wire tU27U11Out;
wire tU27U00Out;
wire tU27U114Out;
wire tU27U112Out;
wire tU27U12Out;
wire tU27U110Out;
wire tU27U18Out;
wire tU27U113Out;
wire tU27U17Out;
wire tU27U19Out;
wire tU27U13Out;
wire tU27U111Out;
wire tU27U16Out;
wire tU27U15Out;
or U27U00(tU27U00Out,tU27U10Out,tU27U11Out,tU27U12Out,tU27U13Out,tU27U14Out,tU27U15Out,tU27U16Out,tU27U17Out,tU27U18Out,tU27U19Out,tU27U110Out,tU27U111Out,tU27U112Out,tU27U113Out,tU27U114Out,tU27U115Out);
and U27U10(tU27U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U27U11(tU27U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U12(tU27U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U27U13(tU27U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U14(tU27U14Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U15(tU27U15Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U16(tU27U16Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U27U17(tU27U17Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U18(tU27U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U27U19(tU27U19Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U110(tU27U110Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U27U111(tU27U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U27U112(tU27U112Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U27U113(tU27U113Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U27U114(tU27U114Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U27U115(tU27U115Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:28====================
wire tU28U120Out;
wire tU28U17Out;
wire tU28U13Out;
wire tU28U110Out;
wire tU28U113Out;
wire tU28U118Out;
wire tU28U18Out;
wire tU28U123Out;
wire tU28U124Out;
wire tU28U114Out;
wire tU28U117Out;
wire tU28U111Out;
wire tU28U115Out;
wire tU28U14Out;
wire tU28U10Out;
wire tU28U116Out;
wire tU28U121Out;
wire tU28U15Out;
wire tU28U122Out;
wire tU28U00Out;
wire tU28U16Out;
wire tU28U112Out;
wire tU28U11Out;
wire tU28U119Out;
wire tU28U12Out;
wire tU28U19Out;
or U28U00(tU28U00Out,tU28U10Out,tU28U11Out,tU28U12Out,tU28U13Out,tU28U14Out,tU28U15Out,tU28U16Out,tU28U17Out,tU28U18Out,tU28U19Out,tU28U110Out,tU28U111Out,tU28U112Out,tU28U113Out,tU28U114Out,tU28U115Out,tU28U116Out,tU28U117Out,tU28U118Out,tU28U119Out,tU28U120Out,tU28U121Out,tU28U122Out,tU28U123Out,tU28U124Out);
and U28U10(tU28U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U28U11(tU28U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U12(tU28U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U13(tU28U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U14(tU28U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U15(tU28U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U16(tU28U16Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U17(tU28U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U18(tU28U18Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U19(tU28U19Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U28U110(tU28U110Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U28U111(tU28U111Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U112(tU28U112Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U113(tU28U113Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U28U114(tU28U114Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U115(tU28U115Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U28U116(tU28U116Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U117(tU28U117Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U28U118(tU28U118Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U28U119(tU28U119Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U28U120(tU28U120Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U28U121(tU28U121Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U28U122(tU28U122Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U28U123(tU28U123Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U28U124(tU28U124Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:29====================
wire tU29U00Out;
wire tU29U110Out;
wire tU29U14Out;
wire tU29U116Out;
wire tU29U112Out;
wire tU29U113Out;
wire tU29U111Out;
wire tU29U115Out;
wire tU29U17Out;
wire tU29U117Out;
wire tU29U118Out;
wire tU29U10Out;
wire tU29U11Out;
wire tU29U114Out;
wire tU29U13Out;
wire tU29U15Out;
wire tU29U12Out;
wire tU29U19Out;
wire tU29U16Out;
wire tU29U18Out;
or U29U00(tU29U00Out,tU29U10Out,tU29U11Out,tU29U12Out,tU29U13Out,tU29U14Out,tU29U15Out,tU29U16Out,tU29U17Out,tU29U18Out,tU29U19Out,tU29U110Out,tU29U111Out,tU29U112Out,tU29U113Out,tU29U114Out,tU29U115Out,tU29U116Out,tU29U117Out,tU29U118Out);
and U29U10(tU29U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U29U11(tU29U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U12(tU29U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U29U13(tU29U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U14(tU29U14Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U15(tU29U15Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U29U16(tU29U16Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U29U17(tU29U17Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U29U18(tU29U18Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U19(tU29U19Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U29U110(tU29U110Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U111(tU29U111Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U112(tU29U112Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U29U113(tU29U113Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U29U114(tU29U114Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U29U115(tU29U115Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U29U116(tU29U116Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U29U117(tU29U117Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U29U118(tU29U118Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:30====================
wire tU30U18Out;
wire tU30U19Out;
wire tU30U116Out;
wire tU30U113Out;
wire tU30U118Out;
wire tU30U111Out;
wire tU30U119Out;
wire tU30U12Out;
wire tU30U120Out;
wire tU30U123Out;
wire tU30U15Out;
wire tU30U11Out;
wire tU30U14Out;
wire tU30U115Out;
wire tU30U00Out;
wire tU30U121Out;
wire tU30U112Out;
wire tU30U16Out;
wire tU30U117Out;
wire tU30U13Out;
wire tU30U17Out;
wire tU30U124Out;
wire tU30U125Out;
wire tU30U126Out;
wire tU30U122Out;
wire tU30U10Out;
wire tU30U110Out;
wire tU30U114Out;
or U30U00(tU30U00Out,tU30U10Out,tU30U11Out,tU30U12Out,tU30U13Out,tU30U14Out,tU30U15Out,tU30U16Out,tU30U17Out,tU30U18Out,tU30U19Out,tU30U110Out,tU30U111Out,tU30U112Out,tU30U113Out,tU30U114Out,tU30U115Out,tU30U116Out,tU30U117Out,tU30U118Out,tU30U119Out,tU30U120Out,tU30U121Out,tU30U122Out,tU30U123Out,tU30U124Out,tU30U125Out,tU30U126Out);
and U30U10(tU30U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U30U11(tU30U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U12(tU30U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U13(tU30U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U14(tU30U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U15(tU30U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U16(tU30U16Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U17(tU30U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U18(tU30U18Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U19(tU30U19Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U30U110(tU30U110Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U30U111(tU30U111Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U30U112(tU30U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U30U113(tU30U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U114(tU30U114Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U115(tU30U115Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U30U116(tU30U116Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U117(tU30U117Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U30U118(tU30U118Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U119(tU30U119Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U30U120(tU30U120Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U30U121(tU30U121Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U30U122(tU30U122Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U30U123(tU30U123Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U30U124(tU30U124Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U30U125(tU30U125Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U30U126(tU30U126Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:31====================
wire tU31U16Out;
wire tU31U18Out;
wire tU31U116Out;
wire tU31U110Out;
wire tU31U11Out;
wire tU31U112Out;
wire tU31U00Out;
wire tU31U114Out;
wire tU31U13Out;
wire tU31U14Out;
wire tU31U17Out;
wire tU31U118Out;
wire tU31U15Out;
wire tU31U12Out;
wire tU31U19Out;
wire tU31U115Out;
wire tU31U111Out;
wire tU31U113Out;
wire tU31U10Out;
wire tU31U117Out;
or U31U00(tU31U00Out,tU31U10Out,tU31U11Out,tU31U12Out,tU31U13Out,tU31U14Out,tU31U15Out,tU31U16Out,tU31U17Out,tU31U18Out,tU31U19Out,tU31U110Out,tU31U111Out,tU31U112Out,tU31U113Out,tU31U114Out,tU31U115Out,tU31U116Out,tU31U117Out,tU31U118Out);
and U31U10(tU31U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U11(tU31U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U12(tU31U12Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U13(tU31U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U14(tU31U14Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U15(tU31U15Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U16(tU31U16Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U17(tU31U17Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U18(tU31U18Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U19(tU31U19Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U31U110(tU31U110Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U111(tU31U111Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U112(tU31U112Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U31U113(tU31U113Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U31U114(tU31U114Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U115(tU31U115Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U31U116(tU31U116Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U31U117(tU31U117Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U31U118(tU31U118Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:32====================
wire tU32U110Out;
wire tU32U12Out;
wire tU32U15Out;
wire tU32U10Out;
wire tU32U19Out;
wire tU32U120Out;
wire tU32U16Out;
wire tU32U111Out;
wire tU32U14Out;
wire tU32U17Out;
wire tU32U00Out;
wire tU32U18Out;
wire tU32U13Out;
wire tU32U118Out;
wire tU32U116Out;
wire tU32U113Out;
wire tU32U119Out;
wire tU32U114Out;
wire tU32U121Out;
wire tU32U117Out;
wire tU32U11Out;
wire tU32U112Out;
wire tU32U115Out;
or U32U00(tU32U00Out,tU32U10Out,tU32U11Out,tU32U12Out,tU32U13Out,tU32U14Out,tU32U15Out,tU32U16Out,tU32U17Out,tU32U18Out,tU32U19Out,tU32U110Out,tU32U111Out,tU32U112Out,tU32U113Out,tU32U114Out,tU32U115Out,tU32U116Out,tU32U117Out,tU32U118Out,tU32U119Out,tU32U120Out,tU32U121Out);
and U32U10(tU32U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U11(tU32U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U12(tU32U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U32U13(tU32U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U32U14(tU32U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U15(tU32U15Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U16(tU32U16Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U32U17(tU32U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U32U18(tU32U18Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U19(tU32U19Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U32U110(tU32U110Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U111(tU32U111Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U112(tU32U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U113(tU32U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U114(tU32U114Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U115(tU32U115Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U32U116(tU32U116Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U117(tU32U117Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U118(tU32U118Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U32U119(tU32U119Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U32U120(tU32U120Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U32U121(tU32U121Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:33====================
wire tU33U17Out;
wire tU33U113Out;
wire tU33U19Out;
wire tU33U00Out;
wire tU33U11Out;
wire tU33U14Out;
wire tU33U112Out;
wire tU33U110Out;
wire tU33U18Out;
wire tU33U10Out;
wire tU33U13Out;
wire tU33U16Out;
wire tU33U15Out;
wire tU33U12Out;
wire tU33U114Out;
wire tU33U111Out;
wire tU33U115Out;
or U33U00(tU33U00Out,tU33U10Out,tU33U11Out,tU33U12Out,tU33U13Out,tU33U14Out,tU33U15Out,tU33U16Out,tU33U17Out,tU33U18Out,tU33U19Out,tU33U110Out,tU33U111Out,tU33U112Out,tU33U113Out,tU33U114Out,tU33U115Out);
and U33U10(tU33U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U11(tU33U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U33U12(tU33U12Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U33U13(tU33U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U14(tU33U14Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U33U15(tU33U15Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U16(tU33U16Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U17(tU33U17Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U18(tU33U18Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U33U19(tU33U19Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U33U110(tU33U110Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U33U111(tU33U111Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U112(tU33U112Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U33U113(tU33U113Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U33U114(tU33U114Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U33U115(tU33U115Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:34====================
wire tU34U126Out;
wire tU34U119Out;
wire tU34U117Out;
wire tU34U18Out;
wire tU34U111Out;
wire tU34U112Out;
wire tU34U116Out;
wire tU34U123Out;
wire tU34U16Out;
wire tU34U13Out;
wire tU34U114Out;
wire tU34U120Out;
wire tU34U125Out;
wire tU34U122Out;
wire tU34U17Out;
wire tU34U127Out;
wire tU34U12Out;
wire tU34U14Out;
wire tU34U00Out;
wire tU34U124Out;
wire tU34U113Out;
wire tU34U115Out;
wire tU34U15Out;
wire tU34U19Out;
wire tU34U11Out;
wire tU34U121Out;
wire tU34U118Out;
wire tU34U10Out;
wire tU34U110Out;
or U34U00(tU34U00Out,tU34U10Out,tU34U11Out,tU34U12Out,tU34U13Out,tU34U14Out,tU34U15Out,tU34U16Out,tU34U17Out,tU34U18Out,tU34U19Out,tU34U110Out,tU34U111Out,tU34U112Out,tU34U113Out,tU34U114Out,tU34U115Out,tU34U116Out,tU34U117Out,tU34U118Out,tU34U119Out,tU34U120Out,tU34U121Out,tU34U122Out,tU34U123Out,tU34U124Out,tU34U125Out,tU34U126Out,tU34U127Out);
and U34U10(tU34U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U11(tU34U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U12(tU34U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U13(tU34U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U14(tU34U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U15(tU34U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U16(tU34U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U17(tU34U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U18(tU34U18Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U19(tU34U19Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U110(tU34U110Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U34U111(tU34U111Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U112(tU34U112Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U113(tU34U113Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U114(tU34U114Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U115(tU34U115Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U116(tU34U116Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U117(tU34U117Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U34U118(tU34U118Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U119(tU34U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U34U120(tU34U120Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U121(tU34U121Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U34U122(tU34U122Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U34U123(tU34U123Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U34U124(tU34U124Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U34U125(tU34U125Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U34U126(tU34U126Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U34U127(tU34U127Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:35====================
wire tU35U120Out;
wire tU35U19Out;
wire tU35U12Out;
wire tU35U16Out;
wire tU35U115Out;
wire tU35U15Out;
wire tU35U118Out;
wire tU35U111Out;
wire tU35U14Out;
wire tU35U00Out;
wire tU35U10Out;
wire tU35U113Out;
wire tU35U117Out;
wire tU35U18Out;
wire tU35U13Out;
wire tU35U114Out;
wire tU35U112Out;
wire tU35U110Out;
wire tU35U116Out;
wire tU35U119Out;
wire tU35U121Out;
wire tU35U11Out;
wire tU35U17Out;
or U35U00(tU35U00Out,tU35U10Out,tU35U11Out,tU35U12Out,tU35U13Out,tU35U14Out,tU35U15Out,tU35U16Out,tU35U17Out,tU35U18Out,tU35U19Out,tU35U110Out,tU35U111Out,tU35U112Out,tU35U113Out,tU35U114Out,tU35U115Out,tU35U116Out,tU35U117Out,tU35U118Out,tU35U119Out,tU35U120Out,tU35U121Out);
and U35U10(tU35U10Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U35U11(tU35U11Out,counter[5],counter[6]);
and U35U12(tU35U12Out,counter[2],counter[4],counter[6]);
and U35U13(tU35U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U35U14(tU35U14Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U35U15(tU35U15Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U35U16(tU35U16Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U35U17(tU35U17Out,counter[2],~counter[4],counter[5]);
and U35U18(tU35U18Out,~counter[1],~counter[3],counter[4],counter[5]);
and U35U19(tU35U19Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U35U110(tU35U110Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U35U111(tU35U111Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U35U112(tU35U112Out,~counter[4],~counter[5],counter[6]);
and U35U113(tU35U113Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U35U114(tU35U114Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U35U115(tU35U115Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U35U116(tU35U116Out,~counter[1],~counter[5],counter[6]);
and U35U117(tU35U117Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U35U118(tU35U118Out,counter[1],~counter[2],counter[4],counter[6]);
and U35U119(tU35U119Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U35U120(tU35U120Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U35U121(tU35U121Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:36====================
wire tU36U10Out;
wire tU36U14Out;
wire tU36U130Out;
wire tU36U111Out;
wire tU36U00Out;
wire tU36U112Out;
wire tU36U118Out;
wire tU36U121Out;
wire tU36U131Out;
wire tU36U124Out;
wire tU36U119Out;
wire tU36U126Out;
wire tU36U113Out;
wire tU36U110Out;
wire tU36U18Out;
wire tU36U123Out;
wire tU36U128Out;
wire tU36U120Out;
wire tU36U17Out;
wire tU36U11Out;
wire tU36U122Out;
wire tU36U15Out;
wire tU36U127Out;
wire tU36U12Out;
wire tU36U16Out;
wire tU36U114Out;
wire tU36U117Out;
wire tU36U19Out;
wire tU36U129Out;
wire tU36U13Out;
wire tU36U115Out;
wire tU36U116Out;
wire tU36U125Out;
or U36U00(tU36U00Out,tU36U10Out,tU36U11Out,tU36U12Out,tU36U13Out,tU36U14Out,tU36U15Out,tU36U16Out,tU36U17Out,tU36U18Out,tU36U19Out,tU36U110Out,tU36U111Out,tU36U112Out,tU36U113Out,tU36U114Out,tU36U115Out,tU36U116Out,tU36U117Out,tU36U118Out,tU36U119Out,tU36U120Out,tU36U121Out,tU36U122Out,tU36U123Out,tU36U124Out,tU36U125Out,tU36U126Out,tU36U127Out,tU36U128Out,tU36U129Out,tU36U130Out,tU36U131Out);
and U36U10(tU36U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U11(tU36U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U12(tU36U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U13(tU36U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U14(tU36U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U15(tU36U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U16(tU36U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U17(tU36U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U18(tU36U18Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U19(tU36U19Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U110(tU36U110Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U36U111(tU36U111Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U112(tU36U112Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U113(tU36U113Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U114(tU36U114Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U115(tU36U115Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U116(tU36U116Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U36U117(tU36U117Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U118(tU36U118Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U36U119(tU36U119Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U120(tU36U120Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U36U121(tU36U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U36U122(tU36U122Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U36U123(tU36U123Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U36U124(tU36U124Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U125(tU36U125Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U36U126(tU36U126Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U36U127(tU36U127Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U36U128(tU36U128Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U36U129(tU36U129Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U36U130(tU36U130Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U36U131(tU36U131Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:37====================
wire tU37U113Out;
wire tU37U00Out;
wire tU37U13Out;
wire tU37U16Out;
wire tU37U18Out;
wire tU37U116Out;
wire tU37U111Out;
wire tU37U112Out;
wire tU37U110Out;
wire tU37U115Out;
wire tU37U19Out;
wire tU37U15Out;
wire tU37U114Out;
wire tU37U12Out;
wire tU37U17Out;
wire tU37U11Out;
wire tU37U10Out;
wire tU37U14Out;
or U37U00(tU37U00Out,tU37U10Out,tU37U11Out,tU37U12Out,tU37U13Out,tU37U14Out,tU37U15Out,tU37U16Out,tU37U17Out,tU37U18Out,tU37U19Out,tU37U110Out,tU37U111Out,tU37U112Out,tU37U113Out,tU37U114Out,tU37U115Out,tU37U116Out);
and U37U10(tU37U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U11(tU37U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U37U12(tU37U12Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U37U13(tU37U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U14(tU37U14Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U15(tU37U15Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U16(tU37U16Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U17(tU37U17Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U37U18(tU37U18Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U37U19(tU37U19Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U37U110(tU37U110Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U37U111(tU37U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U37U112(tU37U112Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U113(tU37U113Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U37U114(tU37U114Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U37U115(tU37U115Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U37U116(tU37U116Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:38====================
wire tU38U122Out;
wire tU38U113Out;
wire tU38U14Out;
wire tU38U117Out;
wire tU38U10Out;
wire tU38U121Out;
wire tU38U18Out;
wire tU38U19Out;
wire tU38U16Out;
wire tU38U123Out;
wire tU38U00Out;
wire tU38U12Out;
wire tU38U110Out;
wire tU38U120Out;
wire tU38U13Out;
wire tU38U116Out;
wire tU38U118Out;
wire tU38U15Out;
wire tU38U115Out;
wire tU38U11Out;
wire tU38U119Out;
wire tU38U17Out;
wire tU38U124Out;
wire tU38U112Out;
wire tU38U114Out;
wire tU38U111Out;
or U38U00(tU38U00Out,tU38U10Out,tU38U11Out,tU38U12Out,tU38U13Out,tU38U14Out,tU38U15Out,tU38U16Out,tU38U17Out,tU38U18Out,tU38U19Out,tU38U110Out,tU38U111Out,tU38U112Out,tU38U113Out,tU38U114Out,tU38U115Out,tU38U116Out,tU38U117Out,tU38U118Out,tU38U119Out,tU38U120Out,tU38U121Out,tU38U122Out,tU38U123Out,tU38U124Out);
and U38U10(tU38U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U11(tU38U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U12(tU38U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U38U13(tU38U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U38U14(tU38U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U15(tU38U15Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U16(tU38U16Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U17(tU38U17Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U18(tU38U18Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U19(tU38U19Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U110(tU38U110Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U111(tU38U111Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U112(tU38U112Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U38U113(tU38U113Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U38U114(tU38U114Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U115(tU38U115Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U38U116(tU38U116Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U38U117(tU38U117Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U118(tU38U118Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U38U119(tU38U119Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U38U120(tU38U120Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U38U121(tU38U121Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U38U122(tU38U122Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U38U123(tU38U123Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U38U124(tU38U124Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:39====================
wire tU39U15Out;
wire tU39U14Out;
wire tU39U11Out;
wire tU39U115Out;
wire tU39U118Out;
wire tU39U117Out;
wire tU39U00Out;
wire tU39U111Out;
wire tU39U18Out;
wire tU39U17Out;
wire tU39U13Out;
wire tU39U114Out;
wire tU39U12Out;
wire tU39U119Out;
wire tU39U110Out;
wire tU39U10Out;
wire tU39U16Out;
wire tU39U112Out;
wire tU39U19Out;
wire tU39U113Out;
wire tU39U116Out;
or U39U00(tU39U00Out,tU39U10Out,tU39U11Out,tU39U12Out,tU39U13Out,tU39U14Out,tU39U15Out,tU39U16Out,tU39U17Out,tU39U18Out,tU39U19Out,tU39U110Out,tU39U111Out,tU39U112Out,tU39U113Out,tU39U114Out,tU39U115Out,tU39U116Out,tU39U117Out,tU39U118Out,tU39U119Out);
and U39U10(tU39U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U11(tU39U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U39U12(tU39U12Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U13(tU39U13Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U39U14(tU39U14Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U15(tU39U15Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U16(tU39U16Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U17(tU39U17Out,~counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U39U18(tU39U18Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U39U19(tU39U19Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U39U110(tU39U110Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U39U111(tU39U111Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U39U112(tU39U112Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U39U113(tU39U113Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U39U114(tU39U114Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U115(tU39U115Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U39U116(tU39U116Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U39U117(tU39U117Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U39U118(tU39U118Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U39U119(tU39U119Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:40====================
wire tU40U10Out;
wire tU40U122Out;
wire tU40U128Out;
wire tU40U12Out;
wire tU40U129Out;
wire tU40U13Out;
wire tU40U133Out;
wire tU40U111Out;
wire tU40U116Out;
wire tU40U11Out;
wire tU40U14Out;
wire tU40U113Out;
wire tU40U118Out;
wire tU40U130Out;
wire tU40U131Out;
wire tU40U127Out;
wire tU40U19Out;
wire tU40U17Out;
wire tU40U112Out;
wire tU40U16Out;
wire tU40U132Out;
wire tU40U00Out;
wire tU40U135Out;
wire tU40U114Out;
wire tU40U134Out;
wire tU40U123Out;
wire tU40U125Out;
wire tU40U110Out;
wire tU40U119Out;
wire tU40U124Out;
wire tU40U115Out;
wire tU40U120Out;
wire tU40U18Out;
wire tU40U15Out;
wire tU40U117Out;
wire tU40U121Out;
wire tU40U126Out;
or U40U00(tU40U00Out,tU40U10Out,tU40U11Out,tU40U12Out,tU40U13Out,tU40U14Out,tU40U15Out,tU40U16Out,tU40U17Out,tU40U18Out,tU40U19Out,tU40U110Out,tU40U111Out,tU40U112Out,tU40U113Out,tU40U114Out,tU40U115Out,tU40U116Out,tU40U117Out,tU40U118Out,tU40U119Out,tU40U120Out,tU40U121Out,tU40U122Out,tU40U123Out,tU40U124Out,tU40U125Out,tU40U126Out,tU40U127Out,tU40U128Out,tU40U129Out,tU40U130Out,tU40U131Out,tU40U132Out,tU40U133Out,tU40U134Out,tU40U135Out);
and U40U10(tU40U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U11(tU40U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U12(tU40U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U40U13(tU40U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U40U14(tU40U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U40U15(tU40U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U16(tU40U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U17(tU40U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U40U18(tU40U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U40U19(tU40U19Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U40U110(tU40U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U111(tU40U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U40U112(tU40U112Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U113(tU40U113Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U114(tU40U114Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U115(tU40U115Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U116(tU40U116Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U40U117(tU40U117Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U40U118(tU40U118Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U119(tU40U119Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U40U120(tU40U120Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U40U121(tU40U121Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U122(tU40U122Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U40U123(tU40U123Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U40U124(tU40U124Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U40U125(tU40U125Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U40U126(tU40U126Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U127(tU40U127Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U40U128(tU40U128Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U40U129(tU40U129Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U40U130(tU40U130Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U40U131(tU40U131Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U40U132(tU40U132Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U40U133(tU40U133Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U40U134(tU40U134Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U40U135(tU40U135Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:41====================
wire tU41U111Out;
wire tU41U122Out;
wire tU41U125Out;
wire tU41U127Out;
wire tU41U124Out;
wire tU41U15Out;
wire tU41U119Out;
wire tU41U00Out;
wire tU41U10Out;
wire tU41U120Out;
wire tU41U110Out;
wire tU41U11Out;
wire tU41U18Out;
wire tU41U121Out;
wire tU41U112Out;
wire tU41U115Out;
wire tU41U117Out;
wire tU41U12Out;
wire tU41U14Out;
wire tU41U16Out;
wire tU41U114Out;
wire tU41U126Out;
wire tU41U19Out;
wire tU41U17Out;
wire tU41U113Out;
wire tU41U13Out;
wire tU41U123Out;
wire tU41U116Out;
wire tU41U118Out;
or U41U00(tU41U00Out,tU41U10Out,tU41U11Out,tU41U12Out,tU41U13Out,tU41U14Out,tU41U15Out,tU41U16Out,tU41U17Out,tU41U18Out,tU41U19Out,tU41U110Out,tU41U111Out,tU41U112Out,tU41U113Out,tU41U114Out,tU41U115Out,tU41U116Out,tU41U117Out,tU41U118Out,tU41U119Out,tU41U120Out,tU41U121Out,tU41U122Out,tU41U123Out,tU41U124Out,tU41U125Out,tU41U126Out,tU41U127Out);
and U41U10(tU41U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U11(tU41U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U41U12(tU41U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U41U13(tU41U13Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U41U14(tU41U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U15(tU41U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U41U16(tU41U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U41U17(tU41U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U41U18(tU41U18Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U41U19(tU41U19Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U41U110(tU41U110Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U111(tU41U111Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U112(tU41U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U113(tU41U113Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U41U114(tU41U114Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U41U115(tU41U115Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U41U116(tU41U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U41U117(tU41U117Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U41U118(tU41U118Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U41U119(tU41U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U41U120(tU41U120Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U41U121(tU41U121Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U122(tU41U122Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U41U123(tU41U123Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U41U124(tU41U124Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U41U125(tU41U125Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U41U126(tU41U126Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U41U127(tU41U127Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:42====================
wire tU42U130Out;
wire tU42U122Out;
wire tU42U123Out;
wire tU42U133Out;
wire tU42U127Out;
wire tU42U15Out;
wire tU42U128Out;
wire tU42U131Out;
wire tU42U115Out;
wire tU42U129Out;
wire tU42U137Out;
wire tU42U10Out;
wire tU42U119Out;
wire tU42U14Out;
wire tU42U13Out;
wire tU42U118Out;
wire tU42U120Out;
wire tU42U16Out;
wire tU42U134Out;
wire tU42U136Out;
wire tU42U110Out;
wire tU42U18Out;
wire tU42U116Out;
wire tU42U00Out;
wire tU42U114Out;
wire tU42U125Out;
wire tU42U112Out;
wire tU42U19Out;
wire tU42U11Out;
wire tU42U12Out;
wire tU42U111Out;
wire tU42U117Out;
wire tU42U135Out;
wire tU42U132Out;
wire tU42U124Out;
wire tU42U126Out;
wire tU42U121Out;
wire tU42U17Out;
wire tU42U113Out;
or U42U00(tU42U00Out,tU42U10Out,tU42U11Out,tU42U12Out,tU42U13Out,tU42U14Out,tU42U15Out,tU42U16Out,tU42U17Out,tU42U18Out,tU42U19Out,tU42U110Out,tU42U111Out,tU42U112Out,tU42U113Out,tU42U114Out,tU42U115Out,tU42U116Out,tU42U117Out,tU42U118Out,tU42U119Out,tU42U120Out,tU42U121Out,tU42U122Out,tU42U123Out,tU42U124Out,tU42U125Out,tU42U126Out,tU42U127Out,tU42U128Out,tU42U129Out,tU42U130Out,tU42U131Out,tU42U132Out,tU42U133Out,tU42U134Out,tU42U135Out,tU42U136Out,tU42U137Out);
and U42U10(tU42U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U11(tU42U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U12(tU42U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U42U13(tU42U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U42U14(tU42U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U42U15(tU42U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U16(tU42U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U17(tU42U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U42U18(tU42U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U42U19(tU42U19Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U42U110(tU42U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U111(tU42U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U42U112(tU42U112Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U42U113(tU42U113Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U114(tU42U114Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U115(tU42U115Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U116(tU42U116Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U117(tU42U117Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U42U118(tU42U118Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U42U119(tU42U119Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U120(tU42U120Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U42U121(tU42U121Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U42U122(tU42U122Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U123(tU42U123Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U42U124(tU42U124Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U42U125(tU42U125Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U42U126(tU42U126Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U42U127(tU42U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U42U128(tU42U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U129(tU42U129Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U42U130(tU42U130Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U42U131(tU42U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U42U132(tU42U132Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U42U133(tU42U133Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U42U134(tU42U134Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U42U135(tU42U135Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U42U136(tU42U136Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U42U137(tU42U137Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:43====================
wire tU43U19Out;
wire tU43U113Out;
wire tU43U15Out;
wire tU43U18Out;
wire tU43U121Out;
wire tU43U111Out;
wire tU43U112Out;
wire tU43U12Out;
wire tU43U115Out;
wire tU43U117Out;
wire tU43U110Out;
wire tU43U17Out;
wire tU43U122Out;
wire tU43U124Out;
wire tU43U00Out;
wire tU43U14Out;
wire tU43U13Out;
wire tU43U16Out;
wire tU43U116Out;
wire tU43U125Out;
wire tU43U123Out;
wire tU43U10Out;
wire tU43U119Out;
wire tU43U118Out;
wire tU43U114Out;
wire tU43U120Out;
wire tU43U11Out;
or U43U00(tU43U00Out,tU43U10Out,tU43U11Out,tU43U12Out,tU43U13Out,tU43U14Out,tU43U15Out,tU43U16Out,tU43U17Out,tU43U18Out,tU43U19Out,tU43U110Out,tU43U111Out,tU43U112Out,tU43U113Out,tU43U114Out,tU43U115Out,tU43U116Out,tU43U117Out,tU43U118Out,tU43U119Out,tU43U120Out,tU43U121Out,tU43U122Out,tU43U123Out,tU43U124Out,tU43U125Out);
and U43U10(tU43U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U11(tU43U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U43U12(tU43U12Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U13(tU43U13Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U43U14(tU43U14Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U43U15(tU43U15Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U16(tU43U16Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U17(tU43U17Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U18(tU43U18Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U43U19(tU43U19Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U43U110(tU43U110Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U43U111(tU43U111Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U43U112(tU43U112Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U43U113(tU43U113Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U43U114(tU43U114Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U43U115(tU43U115Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U43U116(tU43U116Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U43U117(tU43U117Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U43U118(tU43U118Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U43U119(tU43U119Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U120(tU43U120Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U43U121(tU43U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U43U122(tU43U122Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U43U123(tU43U123Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U43U124(tU43U124Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U43U125(tU43U125Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:44====================
wire tU44U124Out;
wire tU44U113Out;
wire tU44U14Out;
wire tU44U110Out;
wire tU44U128Out;
wire tU44U13Out;
wire tU44U10Out;
wire tU44U126Out;
wire tU44U119Out;
wire tU44U131Out;
wire tU44U111Out;
wire tU44U11Out;
wire tU44U112Out;
wire tU44U19Out;
wire tU44U130Out;
wire tU44U18Out;
wire tU44U121Out;
wire tU44U125Out;
wire tU44U00Out;
wire tU44U118Out;
wire tU44U16Out;
wire tU44U129Out;
wire tU44U120Out;
wire tU44U114Out;
wire tU44U12Out;
wire tU44U115Out;
wire tU44U117Out;
wire tU44U122Out;
wire tU44U116Out;
wire tU44U127Out;
wire tU44U15Out;
wire tU44U17Out;
wire tU44U123Out;
or U44U00(tU44U00Out,tU44U10Out,tU44U11Out,tU44U12Out,tU44U13Out,tU44U14Out,tU44U15Out,tU44U16Out,tU44U17Out,tU44U18Out,tU44U19Out,tU44U110Out,tU44U111Out,tU44U112Out,tU44U113Out,tU44U114Out,tU44U115Out,tU44U116Out,tU44U117Out,tU44U118Out,tU44U119Out,tU44U120Out,tU44U121Out,tU44U122Out,tU44U123Out,tU44U124Out,tU44U125Out,tU44U126Out,tU44U127Out,tU44U128Out,tU44U129Out,tU44U130Out,tU44U131Out);
and U44U10(tU44U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U11(tU44U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U12(tU44U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U44U13(tU44U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U14(tU44U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U15(tU44U15Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U44U16(tU44U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U44U17(tU44U17Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U18(tU44U18Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U44U19(tU44U19Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U110(tU44U110Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U111(tU44U111Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U112(tU44U112Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U113(tU44U113Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U44U114(tU44U114Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U115(tU44U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U44U116(tU44U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U44U117(tU44U117Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U118(tU44U118Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U44U119(tU44U119Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U44U120(tU44U120Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U44U121(tU44U121Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U44U122(tU44U122Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U123(tU44U123Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U44U124(tU44U124Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U44U125(tU44U125Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U44U126(tU44U126Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U44U127(tU44U127Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U44U128(tU44U128Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U44U129(tU44U129Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U44U130(tU44U130Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U44U131(tU44U131Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:45====================
wire tU45U114Out;
wire tU45U19Out;
wire tU45U00Out;
wire tU45U13Out;
wire tU45U16Out;
wire tU45U17Out;
wire tU45U111Out;
wire tU45U11Out;
wire tU45U116Out;
wire tU45U112Out;
wire tU45U113Out;
wire tU45U14Out;
wire tU45U10Out;
wire tU45U115Out;
wire tU45U117Out;
wire tU45U15Out;
wire tU45U18Out;
wire tU45U110Out;
wire tU45U12Out;
or U45U00(tU45U00Out,tU45U10Out,tU45U11Out,tU45U12Out,tU45U13Out,tU45U14Out,tU45U15Out,tU45U16Out,tU45U17Out,tU45U18Out,tU45U19Out,tU45U110Out,tU45U111Out,tU45U112Out,tU45U113Out,tU45U114Out,tU45U115Out,tU45U116Out,tU45U117Out);
and U45U10(tU45U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U11(tU45U11Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U12(tU45U12Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U45U13(tU45U13Out,~counter[1],counter[3],~counter[4],counter[5]);
and U45U14(tU45U14Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U15(tU45U15Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U16(tU45U16Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U17(tU45U17Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U45U18(tU45U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U45U19(tU45U19Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U45U110(tU45U110Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U45U111(tU45U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U45U112(tU45U112Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U45U113(tU45U113Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U114(tU45U114Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U45U115(tU45U115Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U45U116(tU45U116Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U45U117(tU45U117Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:46====================
wire tU46U12Out;
wire tU46U18Out;
wire tU46U120Out;
wire tU46U121Out;
wire tU46U136Out;
wire tU46U131Out;
wire tU46U115Out;
wire tU46U11Out;
wire tU46U134Out;
wire tU46U16Out;
wire tU46U14Out;
wire tU46U126Out;
wire tU46U00Out;
wire tU46U128Out;
wire tU46U135Out;
wire tU46U17Out;
wire tU46U139Out;
wire tU46U118Out;
wire tU46U132Out;
wire tU46U15Out;
wire tU46U117Out;
wire tU46U138Out;
wire tU46U124Out;
wire tU46U114Out;
wire tU46U113Out;
wire tU46U116Out;
wire tU46U125Out;
wire tU46U137Out;
wire tU46U129Out;
wire tU46U111Out;
wire tU46U119Out;
wire tU46U19Out;
wire tU46U123Out;
wire tU46U122Out;
wire tU46U133Out;
wire tU46U10Out;
wire tU46U112Out;
wire tU46U130Out;
wire tU46U110Out;
wire tU46U127Out;
wire tU46U13Out;
or U46U00(tU46U00Out,tU46U10Out,tU46U11Out,tU46U12Out,tU46U13Out,tU46U14Out,tU46U15Out,tU46U16Out,tU46U17Out,tU46U18Out,tU46U19Out,tU46U110Out,tU46U111Out,tU46U112Out,tU46U113Out,tU46U114Out,tU46U115Out,tU46U116Out,tU46U117Out,tU46U118Out,tU46U119Out,tU46U120Out,tU46U121Out,tU46U122Out,tU46U123Out,tU46U124Out,tU46U125Out,tU46U126Out,tU46U127Out,tU46U128Out,tU46U129Out,tU46U130Out,tU46U131Out,tU46U132Out,tU46U133Out,tU46U134Out,tU46U135Out,tU46U136Out,tU46U137Out,tU46U138Out,tU46U139Out);
and U46U10(tU46U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U11(tU46U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U12(tU46U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U46U13(tU46U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U46U14(tU46U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U46U15(tU46U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U16(tU46U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U17(tU46U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U46U18(tU46U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U46U19(tU46U19Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U46U110(tU46U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U111(tU46U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U46U112(tU46U112Out,~counter[1],counter[3],~counter[4],counter[5]);
and U46U113(tU46U113Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U46U114(tU46U114Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U115(tU46U115Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U116(tU46U116Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U117(tU46U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U118(tU46U118Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U46U119(tU46U119Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U46U120(tU46U120Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U121(tU46U121Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U46U122(tU46U122Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U46U123(tU46U123Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U46U124(tU46U124Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U125(tU46U125Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U46U126(tU46U126Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U46U127(tU46U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U46U128(tU46U128Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U46U129(tU46U129Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U46U130(tU46U130Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U131(tU46U131Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U46U132(tU46U132Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U46U133(tU46U133Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U46U134(tU46U134Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U46U135(tU46U135Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U46U136(tU46U136Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U46U137(tU46U137Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U46U138(tU46U138Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U46U139(tU46U139Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:47====================
wire tU47U13Out;
wire tU47U122Out;
wire tU47U16Out;
wire tU47U125Out;
wire tU47U10Out;
wire tU47U17Out;
wire tU47U113Out;
wire tU47U00Out;
wire tU47U115Out;
wire tU47U120Out;
wire tU47U12Out;
wire tU47U15Out;
wire tU47U123Out;
wire tU47U11Out;
wire tU47U117Out;
wire tU47U110Out;
wire tU47U18Out;
wire tU47U121Out;
wire tU47U112Out;
wire tU47U116Out;
wire tU47U118Out;
wire tU47U124Out;
wire tU47U111Out;
wire tU47U14Out;
wire tU47U19Out;
wire tU47U114Out;
wire tU47U119Out;
or U47U00(tU47U00Out,tU47U10Out,tU47U11Out,tU47U12Out,tU47U13Out,tU47U14Out,tU47U15Out,tU47U16Out,tU47U17Out,tU47U18Out,tU47U19Out,tU47U110Out,tU47U111Out,tU47U112Out,tU47U113Out,tU47U114Out,tU47U115Out,tU47U116Out,tU47U117Out,tU47U118Out,tU47U119Out,tU47U120Out,tU47U121Out,tU47U122Out,tU47U123Out,tU47U124Out,tU47U125Out);
and U47U10(tU47U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U11(tU47U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U47U12(tU47U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U47U13(tU47U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U14(tU47U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U47U15(tU47U15Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U47U16(tU47U16Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U47U17(tU47U17Out,~counter[1],counter[3],~counter[4],counter[5]);
and U47U18(tU47U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U47U19(tU47U19Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U110(tU47U110Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U111(tU47U111Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U112(tU47U112Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U47U113(tU47U113Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U47U114(tU47U114Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U47U115(tU47U115Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U47U116(tU47U116Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U47U117(tU47U117Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U47U118(tU47U118Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U47U119(tU47U119Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U120(tU47U120Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U47U121(tU47U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U47U122(tU47U122Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U47U123(tU47U123Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U47U124(tU47U124Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U47U125(tU47U125Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:48====================
wire tU48U111Out;
wire tU48U12Out;
wire tU48U14Out;
wire tU48U17Out;
wire tU48U16Out;
wire tU48U110Out;
wire tU48U18Out;
wire tU48U10Out;
wire tU48U113Out;
wire tU48U13Out;
wire tU48U19Out;
wire tU48U15Out;
wire tU48U112Out;
wire tU48U11Out;
wire tU48U00Out;
or U48U00(tU48U00Out,tU48U10Out,tU48U11Out,tU48U12Out,tU48U13Out,tU48U14Out,tU48U15Out,tU48U16Out,tU48U17Out,tU48U18Out,tU48U19Out,tU48U110Out,tU48U111Out,tU48U112Out,tU48U113Out);
and U48U10(tU48U10Out,counter[5],counter[6]);
and U48U11(tU48U11Out,counter[2],counter[4],counter[6]);
and U48U12(tU48U12Out,counter[1],~counter[2],counter[4],counter[5]);
and U48U13(tU48U13Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U48U14(tU48U14Out,counter[0],~counter[2],~counter[3],counter[4],counter[5]);
and U48U15(tU48U15Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U48U16(tU48U16Out,~counter[4],~counter[5],counter[6]);
and U48U17(tU48U17Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U48U18(tU48U18Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U48U19(tU48U19Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U48U110(tU48U110Out,~counter[1],~counter[5],counter[6]);
and U48U111(tU48U111Out,counter[1],~counter[2],counter[4],counter[6]);
and U48U112(tU48U112Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U48U113(tU48U113Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:49====================
wire tU49U115Out;
wire tU49U119Out;
wire tU49U111Out;
wire tU49U117Out;
wire tU49U10Out;
wire tU49U16Out;
wire tU49U13Out;
wire tU49U11Out;
wire tU49U19Out;
wire tU49U14Out;
wire tU49U15Out;
wire tU49U18Out;
wire tU49U118Out;
wire tU49U00Out;
wire tU49U12Out;
wire tU49U120Out;
wire tU49U121Out;
wire tU49U112Out;
wire tU49U110Out;
wire tU49U17Out;
wire tU49U114Out;
wire tU49U113Out;
wire tU49U116Out;
or U49U00(tU49U00Out,tU49U10Out,tU49U11Out,tU49U12Out,tU49U13Out,tU49U14Out,tU49U15Out,tU49U16Out,tU49U17Out,tU49U18Out,tU49U19Out,tU49U110Out,tU49U111Out,tU49U112Out,tU49U113Out,tU49U114Out,tU49U115Out,tU49U116Out,tU49U117Out,tU49U118Out,tU49U119Out,tU49U120Out,tU49U121Out);
and U49U10(tU49U10Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U49U11(tU49U11Out,counter[0],counter[3],counter[4],~counter[5],~counter[6]);
and U49U12(tU49U12Out,~counter[1],counter[3],~counter[4],counter[5]);
and U49U13(tU49U13Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U49U14(tU49U14Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U49U15(tU49U15Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U49U16(tU49U16Out,~counter[1],~counter[2],~counter[3],counter[4],counter[5]);
and U49U17(tU49U17Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U49U18(tU49U18Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U49U19(tU49U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U49U110(tU49U110Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U49U111(tU49U111Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U49U112(tU49U112Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U49U113(tU49U113Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U49U114(tU49U114Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U49U115(tU49U115Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U49U116(tU49U116Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U49U117(tU49U117Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U49U118(tU49U118Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U49U119(tU49U119Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U49U120(tU49U120Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U49U121(tU49U121Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);

//====================Truthtable Variable:50====================
wire tU50U14Out;
wire tU50U13Out;
wire tU50U19Out;
wire tU50U17Out;
wire tU50U116Out;
wire tU50U11Out;
wire tU50U120Out;
wire tU50U122Out;
wire tU50U110Out;
wire tU50U18Out;
wire tU50U114Out;
wire tU50U127Out;
wire tU50U16Out;
wire tU50U125Out;
wire tU50U128Out;
wire tU50U121Out;
wire tU50U119Out;
wire tU50U111Out;
wire tU50U115Out;
wire tU50U113Out;
wire tU50U123Out;
wire tU50U126Out;
wire tU50U12Out;
wire tU50U112Out;
wire tU50U10Out;
wire tU50U117Out;
wire tU50U00Out;
wire tU50U124Out;
wire tU50U118Out;
wire tU50U15Out;
or U50U00(tU50U00Out,tU50U10Out,tU50U11Out,tU50U12Out,tU50U13Out,tU50U14Out,tU50U15Out,tU50U16Out,tU50U17Out,tU50U18Out,tU50U19Out,tU50U110Out,tU50U111Out,tU50U112Out,tU50U113Out,tU50U114Out,tU50U115Out,tU50U116Out,tU50U117Out,tU50U118Out,tU50U119Out,tU50U120Out,tU50U121Out,tU50U122Out,tU50U123Out,tU50U124Out,tU50U125Out,tU50U126Out,tU50U127Out,tU50U128Out);
and U50U10(tU50U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U11(tU50U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U50U12(tU50U12Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U50U13(tU50U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U14(tU50U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U50U15(tU50U15Out,~counter[1],counter[3],~counter[4],counter[5]);
and U50U16(tU50U16Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U50U17(tU50U17Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U50U18(tU50U18Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U19(tU50U19Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U50U110(tU50U110Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U111(tU50U111Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U112(tU50U112Out,~counter[1],~counter[2],~counter[3],counter[4],counter[5]);
and U50U113(tU50U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U50U114(tU50U114Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U50U115(tU50U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U50U116(tU50U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U50U117(tU50U117Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U50U118(tU50U118Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U50U119(tU50U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U50U120(tU50U120Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U50U121(tU50U121Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U122(tU50U122Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U50U123(tU50U123Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U50U124(tU50U124Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U50U125(tU50U125Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U50U126(tU50U126Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U50U127(tU50U127Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U50U128(tU50U128Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:51====================
wire tU51U11Out;
wire tU51U17Out;
wire tU51U18Out;
wire tU51U127Out;
wire tU51U129Out;
wire tU51U111Out;
wire tU51U13Out;
wire tU51U15Out;
wire tU51U120Out;
wire tU51U16Out;
wire tU51U114Out;
wire tU51U128Out;
wire tU51U14Out;
wire tU51U122Out;
wire tU51U121Out;
wire tU51U115Out;
wire tU51U10Out;
wire tU51U123Out;
wire tU51U00Out;
wire tU51U125Out;
wire tU51U117Out;
wire tU51U116Out;
wire tU51U118Out;
wire tU51U110Out;
wire tU51U12Out;
wire tU51U113Out;
wire tU51U119Out;
wire tU51U19Out;
wire tU51U124Out;
wire tU51U112Out;
wire tU51U126Out;
or U51U00(tU51U00Out,tU51U10Out,tU51U11Out,tU51U12Out,tU51U13Out,tU51U14Out,tU51U15Out,tU51U16Out,tU51U17Out,tU51U18Out,tU51U19Out,tU51U110Out,tU51U111Out,tU51U112Out,tU51U113Out,tU51U114Out,tU51U115Out,tU51U116Out,tU51U117Out,tU51U118Out,tU51U119Out,tU51U120Out,tU51U121Out,tU51U122Out,tU51U123Out,tU51U124Out,tU51U125Out,tU51U126Out,tU51U127Out,tU51U128Out,tU51U129Out);
and U51U10(tU51U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U51U11(tU51U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U51U12(tU51U12Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U51U13(tU51U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U51U14(tU51U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U51U15(tU51U15Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U51U16(tU51U16Out,counter[0],~counter[2],~counter[3],counter[4],counter[5]);
and U51U17(tU51U17Out,~counter[1],counter[3],~counter[4],counter[5]);
and U51U18(tU51U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U51U19(tU51U19Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U51U110(tU51U110Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U51U111(tU51U111Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U51U112(tU51U112Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U51U113(tU51U113Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U51U114(tU51U114Out,~counter[1],~counter[2],~counter[3],counter[4],counter[5]);
and U51U115(tU51U115Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U51U116(tU51U116Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U51U117(tU51U117Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U51U118(tU51U118Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U51U119(tU51U119Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U51U120(tU51U120Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U51U121(tU51U121Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U51U122(tU51U122Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U51U123(tU51U123Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U51U124(tU51U124Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U51U125(tU51U125Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U51U126(tU51U126Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U51U127(tU51U127Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U51U128(tU51U128Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U51U129(tU51U129Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);

//====================Truthtable Variable:52====================
wire tU52U13Out;
wire tU52U11Out;
wire tU52U133Out;
wire tU52U129Out;
wire tU52U135Out;
wire tU52U119Out;
wire tU52U18Out;
wire tU52U139Out;
wire tU52U121Out;
wire tU52U140Out;
wire tU52U141Out;
wire tU52U116Out;
wire tU52U142Out;
wire tU52U17Out;
wire tU52U128Out;
wire tU52U143Out;
wire tU52U124Out;
wire tU52U134Out;
wire tU52U127Out;
wire tU52U111Out;
wire tU52U16Out;
wire tU52U10Out;
wire tU52U132Out;
wire tU52U110Out;
wire tU52U15Out;
wire tU52U113Out;
wire tU52U138Out;
wire tU52U117Out;
wire tU52U00Out;
wire tU52U130Out;
wire tU52U118Out;
wire tU52U114Out;
wire tU52U122Out;
wire tU52U12Out;
wire tU52U125Out;
wire tU52U115Out;
wire tU52U14Out;
wire tU52U123Out;
wire tU52U19Out;
wire tU52U112Out;
wire tU52U131Out;
wire tU52U136Out;
wire tU52U120Out;
wire tU52U137Out;
wire tU52U126Out;
or U52U00(tU52U00Out,tU52U10Out,tU52U11Out,tU52U12Out,tU52U13Out,tU52U14Out,tU52U15Out,tU52U16Out,tU52U17Out,tU52U18Out,tU52U19Out,tU52U110Out,tU52U111Out,tU52U112Out,tU52U113Out,tU52U114Out,tU52U115Out,tU52U116Out,tU52U117Out,tU52U118Out,tU52U119Out,tU52U120Out,tU52U121Out,tU52U122Out,tU52U123Out,tU52U124Out,tU52U125Out,tU52U126Out,tU52U127Out,tU52U128Out,tU52U129Out,tU52U130Out,tU52U131Out,tU52U132Out,tU52U133Out,tU52U134Out,tU52U135Out,tU52U136Out,tU52U137Out,tU52U138Out,tU52U139Out,tU52U140Out,tU52U141Out,tU52U142Out,tU52U143Out);
and U52U10(tU52U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U11(tU52U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U12(tU52U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U52U13(tU52U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U52U14(tU52U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U52U15(tU52U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U16(tU52U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U17(tU52U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U52U18(tU52U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U52U19(tU52U19Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U52U110(tU52U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U111(tU52U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U52U112(tU52U112Out,counter[0],~counter[2],~counter[3],counter[4],counter[5]);
and U52U113(tU52U113Out,~counter[1],counter[3],~counter[4],counter[5]);
and U52U114(tU52U114Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U52U115(tU52U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U52U116(tU52U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U117(tU52U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U52U118(tU52U118Out,~counter[0],~counter[1],~counter[3],counter[4],counter[5]);
and U52U119(tU52U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U120(tU52U120Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U121(tU52U121Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U122(tU52U122Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U52U123(tU52U123Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U52U124(tU52U124Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U125(tU52U125Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U52U126(tU52U126Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U52U127(tU52U127Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U52U128(tU52U128Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U129(tU52U129Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U52U130(tU52U130Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U52U131(tU52U131Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U52U132(tU52U132Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U52U133(tU52U133Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U52U134(tU52U134Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U135(tU52U135Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U52U136(tU52U136Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U52U137(tU52U137Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U52U138(tU52U138Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U52U139(tU52U139Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U52U140(tU52U140Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U52U141(tU52U141Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U52U142(tU52U142Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U52U143(tU52U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:53====================
wire tU53U16Out;
wire tU53U111Out;
wire tU53U15Out;
wire tU53U113Out;
wire tU53U112Out;
wire tU53U18Out;
wire tU53U120Out;
wire tU53U10Out;
wire tU53U14Out;
wire tU53U17Out;
wire tU53U128Out;
wire tU53U115Out;
wire tU53U119Out;
wire tU53U131Out;
wire tU53U122Out;
wire tU53U124Out;
wire tU53U110Out;
wire tU53U114Out;
wire tU53U130Out;
wire tU53U126Out;
wire tU53U117Out;
wire tU53U118Out;
wire tU53U19Out;
wire tU53U116Out;
wire tU53U121Out;
wire tU53U00Out;
wire tU53U13Out;
wire tU53U127Out;
wire tU53U125Out;
wire tU53U123Out;
wire tU53U12Out;
wire tU53U11Out;
wire tU53U129Out;
or U53U00(tU53U00Out,tU53U10Out,tU53U11Out,tU53U12Out,tU53U13Out,tU53U14Out,tU53U15Out,tU53U16Out,tU53U17Out,tU53U18Out,tU53U19Out,tU53U110Out,tU53U111Out,tU53U112Out,tU53U113Out,tU53U114Out,tU53U115Out,tU53U116Out,tU53U117Out,tU53U118Out,tU53U119Out,tU53U120Out,tU53U121Out,tU53U122Out,tU53U123Out,tU53U124Out,tU53U125Out,tU53U126Out,tU53U127Out,tU53U128Out,tU53U129Out,tU53U130Out,tU53U131Out);
and U53U10(tU53U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U53U11(tU53U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U53U12(tU53U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U53U13(tU53U13Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U53U14(tU53U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U53U15(tU53U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U53U16(tU53U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U53U17(tU53U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U53U18(tU53U18Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U53U19(tU53U19Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U53U110(tU53U110Out,counter[0],~counter[2],~counter[3],counter[4],counter[5]);
and U53U111(tU53U111Out,~counter[1],counter[3],~counter[4],counter[5]);
and U53U112(tU53U112Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U53U113(tU53U113Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U53U114(tU53U114Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U53U115(tU53U115Out,~counter[1],~counter[3],counter[4],counter[5]);
and U53U116(tU53U116Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U53U117(tU53U117Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U53U118(tU53U118Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U53U119(tU53U119Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U53U120(tU53U120Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U53U121(tU53U121Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U53U122(tU53U122Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U53U123(tU53U123Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U53U124(tU53U124Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U53U125(tU53U125Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U53U126(tU53U126Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U53U127(tU53U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U53U128(tU53U128Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U53U129(tU53U129Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U53U130(tU53U130Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U53U131(tU53U131Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:54====================
wire tU54U116Out;
wire tU54U14Out;
wire tU54U117Out;
wire tU54U126Out;
wire tU54U15Out;
wire tU54U110Out;
wire tU54U18Out;
wire tU54U134Out;
wire tU54U13Out;
wire tU54U137Out;
wire tU54U125Out;
wire tU54U122Out;
wire tU54U19Out;
wire tU54U132Out;
wire tU54U130Out;
wire tU54U123Out;
wire tU54U124Out;
wire tU54U115Out;
wire tU54U00Out;
wire tU54U12Out;
wire tU54U133Out;
wire tU54U112Out;
wire tU54U131Out;
wire tU54U17Out;
wire tU54U119Out;
wire tU54U10Out;
wire tU54U127Out;
wire tU54U135Out;
wire tU54U118Out;
wire tU54U120Out;
wire tU54U129Out;
wire tU54U111Out;
wire tU54U11Out;
wire tU54U121Out;
wire tU54U114Out;
wire tU54U128Out;
wire tU54U136Out;
wire tU54U113Out;
wire tU54U16Out;
or U54U00(tU54U00Out,tU54U10Out,tU54U11Out,tU54U12Out,tU54U13Out,tU54U14Out,tU54U15Out,tU54U16Out,tU54U17Out,tU54U18Out,tU54U19Out,tU54U110Out,tU54U111Out,tU54U112Out,tU54U113Out,tU54U114Out,tU54U115Out,tU54U116Out,tU54U117Out,tU54U118Out,tU54U119Out,tU54U120Out,tU54U121Out,tU54U122Out,tU54U123Out,tU54U124Out,tU54U125Out,tU54U126Out,tU54U127Out,tU54U128Out,tU54U129Out,tU54U130Out,tU54U131Out,tU54U132Out,tU54U133Out,tU54U134Out,tU54U135Out,tU54U136Out,tU54U137Out);
and U54U10(tU54U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U11(tU54U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U54U12(tU54U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U54U13(tU54U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U54U14(tU54U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U54U15(tU54U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U54U16(tU54U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U17(tU54U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U54U18(tU54U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U54U19(tU54U19Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U54U110(tU54U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U54U111(tU54U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U54U112(tU54U112Out,counter[0],~counter[2],~counter[3],counter[4],counter[5]);
and U54U113(tU54U113Out,~counter[1],counter[3],~counter[4],counter[5]);
and U54U114(tU54U114Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U54U115(tU54U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U54U116(tU54U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U117(tU54U117Out,~counter[1],~counter[3],counter[4],counter[5]);
and U54U118(tU54U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U54U119(tU54U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U120(tU54U120Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U121(tU54U121Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U54U122(tU54U122Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U54U123(tU54U123Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U54U124(tU54U124Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U54U125(tU54U125Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U54U126(tU54U126Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U54U127(tU54U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U54U128(tU54U128Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U54U129(tU54U129Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U54U130(tU54U130Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U131(tU54U131Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U54U132(tU54U132Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U54U133(tU54U133Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U54U134(tU54U134Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U54U135(tU54U135Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U54U136(tU54U136Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U54U137(tU54U137Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:55====================
wire tU55U14Out;
wire tU55U118Out;
wire tU55U110Out;
wire tU55U11Out;
wire tU55U121Out;
wire tU55U116Out;
wire tU55U124Out;
wire tU55U119Out;
wire tU55U117Out;
wire tU55U125Out;
wire tU55U16Out;
wire tU55U13Out;
wire tU55U18Out;
wire tU55U126Out;
wire tU55U19Out;
wire tU55U17Out;
wire tU55U123Out;
wire tU55U122Out;
wire tU55U00Out;
wire tU55U115Out;
wire tU55U15Out;
wire tU55U120Out;
wire tU55U113Out;
wire tU55U10Out;
wire tU55U111Out;
wire tU55U112Out;
wire tU55U114Out;
wire tU55U12Out;
or U55U00(tU55U00Out,tU55U10Out,tU55U11Out,tU55U12Out,tU55U13Out,tU55U14Out,tU55U15Out,tU55U16Out,tU55U17Out,tU55U18Out,tU55U19Out,tU55U110Out,tU55U111Out,tU55U112Out,tU55U113Out,tU55U114Out,tU55U115Out,tU55U116Out,tU55U117Out,tU55U118Out,tU55U119Out,tU55U120Out,tU55U121Out,tU55U122Out,tU55U123Out,tU55U124Out,tU55U125Out,tU55U126Out);
and U55U10(tU55U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U55U11(tU55U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U55U12(tU55U12Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U55U13(tU55U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U55U14(tU55U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U55U15(tU55U15Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U55U16(tU55U16Out,~counter[1],counter[3],~counter[4],counter[5]);
and U55U17(tU55U17Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U55U18(tU55U18Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U55U19(tU55U19Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U55U110(tU55U110Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U55U111(tU55U111Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U55U112(tU55U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U55U113(tU55U113Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U55U114(tU55U114Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U55U115(tU55U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U55U116(tU55U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U55U117(tU55U117Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U55U118(tU55U118Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U55U119(tU55U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U55U120(tU55U120Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U55U121(tU55U121Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U55U122(tU55U122Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U55U123(tU55U123Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U55U124(tU55U124Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U55U125(tU55U125Out,~counter[3],counter[4],counter[5]);
and U55U126(tU55U126Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);

//====================Truthtable Variable:56====================
wire tU56U127Out;
wire tU56U126Out;
wire tU56U117Out;
wire tU56U111Out;
wire tU56U122Out;
wire tU56U115Out;
wire tU56U116Out;
wire tU56U123Out;
wire tU56U112Out;
wire tU56U10Out;
wire tU56U15Out;
wire tU56U118Out;
wire tU56U120Out;
wire tU56U125Out;
wire tU56U14Out;
wire tU56U16Out;
wire tU56U113Out;
wire tU56U119Out;
wire tU56U11Out;
wire tU56U17Out;
wire tU56U00Out;
wire tU56U124Out;
wire tU56U18Out;
wire tU56U121Out;
wire tU56U13Out;
wire tU56U110Out;
wire tU56U19Out;
wire tU56U12Out;
wire tU56U114Out;
or U56U00(tU56U00Out,tU56U10Out,tU56U11Out,tU56U12Out,tU56U13Out,tU56U14Out,tU56U15Out,tU56U16Out,tU56U17Out,tU56U18Out,tU56U19Out,tU56U110Out,tU56U111Out,tU56U112Out,tU56U113Out,tU56U114Out,tU56U115Out,tU56U116Out,tU56U117Out,tU56U118Out,tU56U119Out,tU56U120Out,tU56U121Out,tU56U122Out,tU56U123Out,tU56U124Out,tU56U125Out,tU56U126Out,tU56U127Out);
and U56U10(tU56U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U56U11(tU56U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U56U12(tU56U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U56U13(tU56U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U56U14(tU56U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U56U15(tU56U15Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U56U16(tU56U16Out,~counter[0],~counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U56U17(tU56U17Out,~counter[1],counter[3],~counter[4],counter[5]);
and U56U18(tU56U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U56U19(tU56U19Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U56U110(tU56U110Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U56U111(tU56U111Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U56U112(tU56U112Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U56U113(tU56U113Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U56U114(tU56U114Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U56U115(tU56U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U56U116(tU56U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U56U117(tU56U117Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U56U118(tU56U118Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U56U119(tU56U119Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U56U120(tU56U120Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U56U121(tU56U121Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U56U122(tU56U122Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U56U123(tU56U123Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U56U124(tU56U124Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U56U125(tU56U125Out,~counter[3],counter[4],counter[5]);
and U56U126(tU56U126Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U56U127(tU56U127Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:57====================
wire tU57U14Out;
wire tU57U19Out;
wire tU57U112Out;
wire tU57U00Out;
wire tU57U113Out;
wire tU57U115Out;
wire tU57U110Out;
wire tU57U18Out;
wire tU57U10Out;
wire tU57U12Out;
wire tU57U117Out;
wire tU57U13Out;
wire tU57U114Out;
wire tU57U17Out;
wire tU57U16Out;
wire tU57U11Out;
wire tU57U116Out;
wire tU57U15Out;
wire tU57U111Out;
or U57U00(tU57U00Out,tU57U10Out,tU57U11Out,tU57U12Out,tU57U13Out,tU57U14Out,tU57U15Out,tU57U16Out,tU57U17Out,tU57U18Out,tU57U19Out,tU57U110Out,tU57U111Out,tU57U112Out,tU57U113Out,tU57U114Out,tU57U115Out,tU57U116Out,tU57U117Out);
and U57U10(tU57U10Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U57U11(tU57U11Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U57U12(tU57U12Out,~counter[1],counter[3],~counter[4],counter[5]);
and U57U13(tU57U13Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U57U14(tU57U14Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U57U15(tU57U15Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U57U16(tU57U16Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U57U17(tU57U17Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U57U18(tU57U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U57U19(tU57U19Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U57U110(tU57U110Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U57U111(tU57U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U57U112(tU57U112Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U57U113(tU57U113Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U57U114(tU57U114Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U57U115(tU57U115Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U57U116(tU57U116Out,~counter[3],counter[4],counter[5]);
and U57U117(tU57U117Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);

//====================Truthtable Variable:58====================
wire tU58U12Out;
wire tU58U115Out;
wire tU58U130Out;
wire tU58U138Out;
wire tU58U11Out;
wire tU58U135Out;
wire tU58U14Out;
wire tU58U124Out;
wire tU58U125Out;
wire tU58U132Out;
wire tU58U141Out;
wire tU58U143Out;
wire tU58U17Out;
wire tU58U18Out;
wire tU58U15Out;
wire tU58U117Out;
wire tU58U128Out;
wire tU58U119Out;
wire tU58U10Out;
wire tU58U110Out;
wire tU58U122Out;
wire tU58U19Out;
wire tU58U116Out;
wire tU58U13Out;
wire tU58U127Out;
wire tU58U131Out;
wire tU58U121Out;
wire tU58U140Out;
wire tU58U129Out;
wire tU58U16Out;
wire tU58U133Out;
wire tU58U112Out;
wire tU58U136Out;
wire tU58U113Out;
wire tU58U126Out;
wire tU58U120Out;
wire tU58U134Out;
wire tU58U123Out;
wire tU58U118Out;
wire tU58U137Out;
wire tU58U142Out;
wire tU58U139Out;
wire tU58U00Out;
wire tU58U111Out;
wire tU58U114Out;
or U58U00(tU58U00Out,tU58U10Out,tU58U11Out,tU58U12Out,tU58U13Out,tU58U14Out,tU58U15Out,tU58U16Out,tU58U17Out,tU58U18Out,tU58U19Out,tU58U110Out,tU58U111Out,tU58U112Out,tU58U113Out,tU58U114Out,tU58U115Out,tU58U116Out,tU58U117Out,tU58U118Out,tU58U119Out,tU58U120Out,tU58U121Out,tU58U122Out,tU58U123Out,tU58U124Out,tU58U125Out,tU58U126Out,tU58U127Out,tU58U128Out,tU58U129Out,tU58U130Out,tU58U131Out,tU58U132Out,tU58U133Out,tU58U134Out,tU58U135Out,tU58U136Out,tU58U137Out,tU58U138Out,tU58U139Out,tU58U140Out,tU58U141Out,tU58U142Out,tU58U143Out);
and U58U10(tU58U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U58U11(tU58U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U58U12(tU58U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U58U13(tU58U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U58U14(tU58U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U58U15(tU58U15Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U58U16(tU58U16Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U58U17(tU58U17Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U58U18(tU58U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U58U19(tU58U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U58U110(tU58U110Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U58U111(tU58U111Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U58U112(tU58U112Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U58U113(tU58U113Out,~counter[1],counter[3],~counter[4],counter[5]);
and U58U114(tU58U114Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U58U115(tU58U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U58U116(tU58U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U58U117(tU58U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U58U118(tU58U118Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U58U119(tU58U119Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U58U120(tU58U120Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U58U121(tU58U121Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U58U122(tU58U122Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U58U123(tU58U123Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U58U124(tU58U124Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U58U125(tU58U125Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U58U126(tU58U126Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U58U127(tU58U127Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U58U128(tU58U128Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U58U129(tU58U129Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U58U130(tU58U130Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U58U131(tU58U131Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U58U132(tU58U132Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U58U133(tU58U133Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U58U134(tU58U134Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U58U135(tU58U135Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U58U136(tU58U136Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U58U137(tU58U137Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U58U138(tU58U138Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U58U139(tU58U139Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U58U140(tU58U140Out,~counter[3],counter[4],counter[5]);
and U58U141(tU58U141Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U58U142(tU58U142Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U58U143(tU58U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:59====================
wire tU59U00Out;
wire tU59U118Out;
wire tU59U16Out;
wire tU59U123Out;
wire tU59U13Out;
wire tU59U121Out;
wire tU59U112Out;
wire tU59U116Out;
wire tU59U122Out;
wire tU59U111Out;
wire tU59U11Out;
wire tU59U18Out;
wire tU59U17Out;
wire tU59U15Out;
wire tU59U113Out;
wire tU59U117Out;
wire tU59U19Out;
wire tU59U124Out;
wire tU59U10Out;
wire tU59U120Out;
wire tU59U115Out;
wire tU59U110Out;
wire tU59U114Out;
wire tU59U12Out;
wire tU59U125Out;
wire tU59U119Out;
wire tU59U14Out;
wire tU59U126Out;
or U59U00(tU59U00Out,tU59U10Out,tU59U11Out,tU59U12Out,tU59U13Out,tU59U14Out,tU59U15Out,tU59U16Out,tU59U17Out,tU59U18Out,tU59U19Out,tU59U110Out,tU59U111Out,tU59U112Out,tU59U113Out,tU59U114Out,tU59U115Out,tU59U116Out,tU59U117Out,tU59U118Out,tU59U119Out,tU59U120Out,tU59U121Out,tU59U122Out,tU59U123Out,tU59U124Out,tU59U125Out,tU59U126Out);
and U59U10(tU59U10Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U59U11(tU59U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U59U12(tU59U12Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U59U13(tU59U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U59U14(tU59U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U59U15(tU59U15Out,counter[1],~counter[2],counter[4],counter[5]);
and U59U16(tU59U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U59U17(tU59U17Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U59U18(tU59U18Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U59U19(tU59U19Out,~counter[1],counter[3],~counter[4],counter[5]);
and U59U110(tU59U110Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U59U111(tU59U111Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U59U112(tU59U112Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U59U113(tU59U113Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U59U114(tU59U114Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U59U115(tU59U115Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U59U116(tU59U116Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U59U117(tU59U117Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U59U118(tU59U118Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U59U119(tU59U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U59U120(tU59U120Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U59U121(tU59U121Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U59U122(tU59U122Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U59U123(tU59U123Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U59U124(tU59U124Out,~counter[3],counter[4],counter[5]);
and U59U125(tU59U125Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U59U126(tU59U126Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:60====================
wire tU60U117Out;
wire tU60U00Out;
wire tU60U115Out;
wire tU60U19Out;
wire tU60U14Out;
wire tU60U110Out;
wire tU60U141Out;
wire tU60U16Out;
wire tU60U116Out;
wire tU60U123Out;
wire tU60U125Out;
wire tU60U127Out;
wire tU60U129Out;
wire tU60U17Out;
wire tU60U143Out;
wire tU60U122Out;
wire tU60U112Out;
wire tU60U130Out;
wire tU60U134Out;
wire tU60U133Out;
wire tU60U126Out;
wire tU60U18Out;
wire tU60U136Out;
wire tU60U119Out;
wire tU60U140Out;
wire tU60U12Out;
wire tU60U13Out;
wire tU60U111Out;
wire tU60U145Out;
wire tU60U114Out;
wire tU60U15Out;
wire tU60U142Out;
wire tU60U11Out;
wire tU60U139Out;
wire tU60U128Out;
wire tU60U138Out;
wire tU60U144Out;
wire tU60U120Out;
wire tU60U118Out;
wire tU60U10Out;
wire tU60U124Out;
wire tU60U132Out;
wire tU60U137Out;
wire tU60U113Out;
wire tU60U121Out;
wire tU60U135Out;
wire tU60U131Out;
or U60U00(tU60U00Out,tU60U10Out,tU60U11Out,tU60U12Out,tU60U13Out,tU60U14Out,tU60U15Out,tU60U16Out,tU60U17Out,tU60U18Out,tU60U19Out,tU60U110Out,tU60U111Out,tU60U112Out,tU60U113Out,tU60U114Out,tU60U115Out,tU60U116Out,tU60U117Out,tU60U118Out,tU60U119Out,tU60U120Out,tU60U121Out,tU60U122Out,tU60U123Out,tU60U124Out,tU60U125Out,tU60U126Out,tU60U127Out,tU60U128Out,tU60U129Out,tU60U130Out,tU60U131Out,tU60U132Out,tU60U133Out,tU60U134Out,tU60U135Out,tU60U136Out,tU60U137Out,tU60U138Out,tU60U139Out,tU60U140Out,tU60U141Out,tU60U142Out,tU60U143Out,tU60U144Out,tU60U145Out);
and U60U10(tU60U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U60U11(tU60U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U60U12(tU60U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U60U13(tU60U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U60U14(tU60U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U60U15(tU60U15Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U60U16(tU60U16Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U60U17(tU60U17Out,~counter[0],~counter[1],counter[3],counter[5]);
and U60U18(tU60U18Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U60U19(tU60U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U60U110(tU60U110Out,counter[1],~counter[2],counter[4],counter[5]);
and U60U111(tU60U111Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U60U112(tU60U112Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U60U113(tU60U113Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U60U114(tU60U114Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U60U115(tU60U115Out,~counter[1],counter[3],~counter[4],counter[5]);
and U60U116(tU60U116Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U60U117(tU60U117Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U60U118(tU60U118Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U60U119(tU60U119Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U60U120(tU60U120Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U60U121(tU60U121Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U60U122(tU60U122Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U60U123(tU60U123Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U60U124(tU60U124Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U60U125(tU60U125Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U60U126(tU60U126Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U60U127(tU60U127Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U60U128(tU60U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U60U129(tU60U129Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U60U130(tU60U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U60U131(tU60U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U60U132(tU60U132Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U60U133(tU60U133Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U60U134(tU60U134Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U60U135(tU60U135Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U60U136(tU60U136Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U60U137(tU60U137Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U60U138(tU60U138Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U60U139(tU60U139Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U60U140(tU60U140Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U60U141(tU60U141Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U60U142(tU60U142Out,~counter[3],counter[4],counter[5]);
and U60U143(tU60U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U60U144(tU60U144Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U60U145(tU60U145Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:61====================
wire tU61U114Out;
wire tU61U14Out;
wire tU61U16Out;
wire tU61U00Out;
wire tU61U111Out;
wire tU61U11Out;
wire tU61U12Out;
wire tU61U118Out;
wire tU61U15Out;
wire tU61U112Out;
wire tU61U113Out;
wire tU61U110Out;
wire tU61U19Out;
wire tU61U116Out;
wire tU61U117Out;
wire tU61U17Out;
wire tU61U13Out;
wire tU61U115Out;
wire tU61U18Out;
wire tU61U10Out;
or U61U00(tU61U00Out,tU61U10Out,tU61U11Out,tU61U12Out,tU61U13Out,tU61U14Out,tU61U15Out,tU61U16Out,tU61U17Out,tU61U18Out,tU61U19Out,tU61U110Out,tU61U111Out,tU61U112Out,tU61U113Out,tU61U114Out,tU61U115Out,tU61U116Out,tU61U117Out,tU61U118Out);
and U61U10(tU61U10Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U61U11(tU61U11Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U61U12(tU61U12Out,counter[1],~counter[2],counter[4],counter[5]);
and U61U13(tU61U13Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U61U14(tU61U14Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U61U15(tU61U15Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U61U16(tU61U16Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U61U17(tU61U17Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U61U18(tU61U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U61U19(tU61U19Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U61U110(tU61U110Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U61U111(tU61U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U61U112(tU61U112Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U61U113(tU61U113Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U61U114(tU61U114Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U61U115(tU61U115Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U61U116(tU61U116Out,~counter[3],counter[4],counter[5]);
and U61U117(tU61U117Out,~counter[1],counter[2],counter[3],counter[5]);
and U61U118(tU61U118Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);

//====================Truthtable Variable:62====================
wire tU62U119Out;
wire tU62U14Out;
wire tU62U128Out;
wire tU62U123Out;
wire tU62U112Out;
wire tU62U00Out;
wire tU62U126Out;
wire tU62U15Out;
wire tU62U115Out;
wire tU62U124Out;
wire tU62U110Out;
wire tU62U121Out;
wire tU62U117Out;
wire tU62U18Out;
wire tU62U19Out;
wire tU62U11Out;
wire tU62U122Out;
wire tU62U127Out;
wire tU62U113Out;
wire tU62U16Out;
wire tU62U111Out;
wire tU62U17Out;
wire tU62U125Out;
wire tU62U13Out;
wire tU62U118Out;
wire tU62U116Out;
wire tU62U12Out;
wire tU62U10Out;
wire tU62U114Out;
wire tU62U129Out;
wire tU62U120Out;
or U62U00(tU62U00Out,tU62U10Out,tU62U11Out,tU62U12Out,tU62U13Out,tU62U14Out,tU62U15Out,tU62U16Out,tU62U17Out,tU62U18Out,tU62U19Out,tU62U110Out,tU62U111Out,tU62U112Out,tU62U113Out,tU62U114Out,tU62U115Out,tU62U116Out,tU62U117Out,tU62U118Out,tU62U119Out,tU62U120Out,tU62U121Out,tU62U122Out,tU62U123Out,tU62U124Out,tU62U125Out,tU62U126Out,tU62U127Out,tU62U128Out,tU62U129Out);
and U62U10(tU62U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U62U11(tU62U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U62U12(tU62U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U62U13(tU62U13Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U62U14(tU62U14Out,counter[1],~counter[2],counter[4],counter[5]);
and U62U15(tU62U15Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U62U16(tU62U16Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U62U17(tU62U17Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U62U18(tU62U18Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U62U19(tU62U19Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U62U110(tU62U110Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U62U111(tU62U111Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U62U112(tU62U112Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U62U113(tU62U113Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U62U114(tU62U114Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U62U115(tU62U115Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U62U116(tU62U116Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U62U117(tU62U117Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U62U118(tU62U118Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U62U119(tU62U119Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U62U120(tU62U120Out,~counter[0],counter[2],counter[3],counter[5]);
and U62U121(tU62U121Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U62U122(tU62U122Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U62U123(tU62U123Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U62U124(tU62U124Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U62U125(tU62U125Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U62U126(tU62U126Out,~counter[3],counter[4],counter[5]);
and U62U127(tU62U127Out,~counter[1],counter[2],counter[3],counter[5]);
and U62U128(tU62U128Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U62U129(tU62U129Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);

//====================Truthtable Variable:63====================
wire tU63U113Out;
wire tU63U110Out;
wire tU63U116Out;
wire tU63U118Out;
wire tU63U119Out;
wire tU63U121Out;
wire tU63U120Out;
wire tU63U123Out;
wire tU63U112Out;
wire tU63U12Out;
wire tU63U00Out;
wire tU63U115Out;
wire tU63U15Out;
wire tU63U18Out;
wire tU63U13Out;
wire tU63U17Out;
wire tU63U19Out;
wire tU63U122Out;
wire tU63U14Out;
wire tU63U10Out;
wire tU63U114Out;
wire tU63U16Out;
wire tU63U117Out;
wire tU63U111Out;
wire tU63U11Out;
or U63U00(tU63U00Out,tU63U10Out,tU63U11Out,tU63U12Out,tU63U13Out,tU63U14Out,tU63U15Out,tU63U16Out,tU63U17Out,tU63U18Out,tU63U19Out,tU63U110Out,tU63U111Out,tU63U112Out,tU63U113Out,tU63U114Out,tU63U115Out,tU63U116Out,tU63U117Out,tU63U118Out,tU63U119Out,tU63U120Out,tU63U121Out,tU63U122Out,tU63U123Out);
and U63U10(tU63U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U11(tU63U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U12(tU63U12Out,counter[5],counter[6]);
and U63U13(tU63U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U14(tU63U14Out,counter[2],counter[4],counter[6]);
and U63U15(tU63U15Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U16(tU63U16Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U17(tU63U17Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U18(tU63U18Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U19(tU63U19Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U110(tU63U110Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U111(tU63U111Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U63U112(tU63U112Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U113(tU63U113Out,~counter[4],~counter[5],counter[6]);
and U63U114(tU63U114Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U115(tU63U115Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U63U116(tU63U116Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U63U117(tU63U117Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U118(tU63U118Out,~counter[1],~counter[5],counter[6]);
and U63U119(tU63U119Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U63U120(tU63U120Out,counter[1],~counter[2],counter[4],counter[6]);
and U63U121(tU63U121Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U63U122(tU63U122Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U63U123(tU63U123Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:64====================
wire tU64U13Out;
wire tU64U135Out;
wire tU64U17Out;
wire tU64U15Out;
wire tU64U116Out;
wire tU64U121Out;
wire tU64U133Out;
wire tU64U138Out;
wire tU64U113Out;
wire tU64U12Out;
wire tU64U132Out;
wire tU64U18Out;
wire tU64U122Out;
wire tU64U131Out;
wire tU64U11Out;
wire tU64U16Out;
wire tU64U110Out;
wire tU64U118Out;
wire tU64U10Out;
wire tU64U127Out;
wire tU64U136Out;
wire tU64U115Out;
wire tU64U134Out;
wire tU64U120Out;
wire tU64U140Out;
wire tU64U137Out;
wire tU64U119Out;
wire tU64U129Out;
wire tU64U00Out;
wire tU64U126Out;
wire tU64U114Out;
wire tU64U19Out;
wire tU64U111Out;
wire tU64U14Out;
wire tU64U123Out;
wire tU64U130Out;
wire tU64U117Out;
wire tU64U124Out;
wire tU64U125Out;
wire tU64U128Out;
wire tU64U139Out;
wire tU64U112Out;
or U64U00(tU64U00Out,tU64U10Out,tU64U11Out,tU64U12Out,tU64U13Out,tU64U14Out,tU64U15Out,tU64U16Out,tU64U17Out,tU64U18Out,tU64U19Out,tU64U110Out,tU64U111Out,tU64U112Out,tU64U113Out,tU64U114Out,tU64U115Out,tU64U116Out,tU64U117Out,tU64U118Out,tU64U119Out,tU64U120Out,tU64U121Out,tU64U122Out,tU64U123Out,tU64U124Out,tU64U125Out,tU64U126Out,tU64U127Out,tU64U128Out,tU64U129Out,tU64U130Out,tU64U131Out,tU64U132Out,tU64U133Out,tU64U134Out,tU64U135Out,tU64U136Out,tU64U137Out,tU64U138Out,tU64U139Out,tU64U140Out);
and U64U10(tU64U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U64U11(tU64U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U64U12(tU64U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U64U13(tU64U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U64U14(tU64U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U64U15(tU64U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U64U16(tU64U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U64U17(tU64U17Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U64U18(tU64U18Out,counter[1],~counter[2],counter[4],counter[5]);
and U64U19(tU64U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U64U110(tU64U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U64U111(tU64U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U64U112(tU64U112Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U64U113(tU64U113Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U64U114(tU64U114Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U64U115(tU64U115Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U64U116(tU64U116Out,~counter[1],~counter[3],counter[4],counter[5]);
and U64U117(tU64U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U64U118(tU64U118Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U64U119(tU64U119Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U64U120(tU64U120Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U64U121(tU64U121Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U64U122(tU64U122Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U64U123(tU64U123Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U64U124(tU64U124Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U64U125(tU64U125Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U64U126(tU64U126Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U64U127(tU64U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U64U128(tU64U128Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U64U129(tU64U129Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U64U130(tU64U130Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U64U131(tU64U131Out,~counter[0],counter[2],counter[3],counter[5]);
and U64U132(tU64U132Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U64U133(tU64U133Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U64U134(tU64U134Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U64U135(tU64U135Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U64U136(tU64U136Out,~counter[1],counter[2],counter[3],counter[5]);
and U64U137(tU64U137Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U64U138(tU64U138Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U64U139(tU64U139Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U64U140(tU64U140Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:65====================
wire tU65U113Out;
wire tU65U128Out;
wire tU65U118Out;
wire tU65U110Out;
wire tU65U16Out;
wire tU65U130Out;
wire tU65U121Out;
wire tU65U129Out;
wire tU65U111Out;
wire tU65U117Out;
wire tU65U125Out;
wire tU65U17Out;
wire tU65U12Out;
wire tU65U114Out;
wire tU65U116Out;
wire tU65U120Out;
wire tU65U122Out;
wire tU65U115Out;
wire tU65U10Out;
wire tU65U11Out;
wire tU65U18Out;
wire tU65U119Out;
wire tU65U131Out;
wire tU65U132Out;
wire tU65U127Out;
wire tU65U00Out;
wire tU65U15Out;
wire tU65U13Out;
wire tU65U124Out;
wire tU65U126Out;
wire tU65U19Out;
wire tU65U112Out;
wire tU65U14Out;
wire tU65U123Out;
or U65U00(tU65U00Out,tU65U10Out,tU65U11Out,tU65U12Out,tU65U13Out,tU65U14Out,tU65U15Out,tU65U16Out,tU65U17Out,tU65U18Out,tU65U19Out,tU65U110Out,tU65U111Out,tU65U112Out,tU65U113Out,tU65U114Out,tU65U115Out,tU65U116Out,tU65U117Out,tU65U118Out,tU65U119Out,tU65U120Out,tU65U121Out,tU65U122Out,tU65U123Out,tU65U124Out,tU65U125Out,tU65U126Out,tU65U127Out,tU65U128Out,tU65U129Out,tU65U130Out,tU65U131Out,tU65U132Out);
and U65U10(tU65U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U65U11(tU65U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U65U12(tU65U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U65U13(tU65U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U65U14(tU65U14Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U65U15(tU65U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U65U16(tU65U16Out,counter[1],~counter[2],counter[4],counter[5]);
and U65U17(tU65U17Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U65U18(tU65U18Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U65U19(tU65U19Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U65U110(tU65U110Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U65U111(tU65U111Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U65U112(tU65U112Out,~counter[1],~counter[3],counter[4],counter[5]);
and U65U113(tU65U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U65U114(tU65U114Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U65U115(tU65U115Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U65U116(tU65U116Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U65U117(tU65U117Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U65U118(tU65U118Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U65U119(tU65U119Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U65U120(tU65U120Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U65U121(tU65U121Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U65U122(tU65U122Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U65U123(tU65U123Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U65U124(tU65U124Out,~counter[0],counter[2],counter[3],counter[5]);
and U65U125(tU65U125Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U65U126(tU65U126Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U65U127(tU65U127Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U65U128(tU65U128Out,~counter[1],counter[2],counter[3],counter[5]);
and U65U129(tU65U129Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U65U130(tU65U130Out,~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U65U131(tU65U131Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U65U132(tU65U132Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:66====================
wire tU66U140Out;
wire tU66U17Out;
wire tU66U133Out;
wire tU66U14Out;
wire tU66U11Out;
wire tU66U137Out;
wire tU66U111Out;
wire tU66U13Out;
wire tU66U120Out;
wire tU66U142Out;
wire tU66U146Out;
wire tU66U15Out;
wire tU66U115Out;
wire tU66U138Out;
wire tU66U141Out;
wire tU66U130Out;
wire tU66U145Out;
wire tU66U124Out;
wire tU66U12Out;
wire tU66U147Out;
wire tU66U116Out;
wire tU66U125Out;
wire tU66U129Out;
wire tU66U19Out;
wire tU66U136Out;
wire tU66U143Out;
wire tU66U10Out;
wire tU66U134Out;
wire tU66U119Out;
wire tU66U114Out;
wire tU66U128Out;
wire tU66U110Out;
wire tU66U131Out;
wire tU66U132Out;
wire tU66U148Out;
wire tU66U18Out;
wire tU66U112Out;
wire tU66U16Out;
wire tU66U118Out;
wire tU66U113Out;
wire tU66U123Out;
wire tU66U126Out;
wire tU66U127Out;
wire tU66U144Out;
wire tU66U117Out;
wire tU66U121Out;
wire tU66U135Out;
wire tU66U139Out;
wire tU66U00Out;
wire tU66U122Out;
or U66U00(tU66U00Out,tU66U10Out,tU66U11Out,tU66U12Out,tU66U13Out,tU66U14Out,tU66U15Out,tU66U16Out,tU66U17Out,tU66U18Out,tU66U19Out,tU66U110Out,tU66U111Out,tU66U112Out,tU66U113Out,tU66U114Out,tU66U115Out,tU66U116Out,tU66U117Out,tU66U118Out,tU66U119Out,tU66U120Out,tU66U121Out,tU66U122Out,tU66U123Out,tU66U124Out,tU66U125Out,tU66U126Out,tU66U127Out,tU66U128Out,tU66U129Out,tU66U130Out,tU66U131Out,tU66U132Out,tU66U133Out,tU66U134Out,tU66U135Out,tU66U136Out,tU66U137Out,tU66U138Out,tU66U139Out,tU66U140Out,tU66U141Out,tU66U142Out,tU66U143Out,tU66U144Out,tU66U145Out,tU66U146Out,tU66U147Out,tU66U148Out);
and U66U10(tU66U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U66U11(tU66U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U66U12(tU66U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U66U13(tU66U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U66U14(tU66U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U66U15(tU66U15Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U66U16(tU66U16Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U66U17(tU66U17Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U66U18(tU66U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U66U19(tU66U19Out,counter[1],~counter[2],counter[4],counter[5]);
and U66U110(tU66U110Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U66U111(tU66U111Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U66U112(tU66U112Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U66U113(tU66U113Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U66U114(tU66U114Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U66U115(tU66U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U66U116(tU66U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U66U117(tU66U117Out,~counter[1],~counter[3],counter[4],counter[5]);
and U66U118(tU66U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U66U119(tU66U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U66U120(tU66U120Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U66U121(tU66U121Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U66U122(tU66U122Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U66U123(tU66U123Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U66U124(tU66U124Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U66U125(tU66U125Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U66U126(tU66U126Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U66U127(tU66U127Out,~counter[0],~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U66U128(tU66U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U66U129(tU66U129Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U66U130(tU66U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U66U131(tU66U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U66U132(tU66U132Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U66U133(tU66U133Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U66U134(tU66U134Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U66U135(tU66U135Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U66U136(tU66U136Out,~counter[0],counter[2],counter[3],counter[5]);
and U66U137(tU66U137Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U66U138(tU66U138Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U66U139(tU66U139Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U66U140(tU66U140Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U66U141(tU66U141Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U66U142(tU66U142Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U66U143(tU66U143Out,~counter[1],counter[2],counter[3],counter[5]);
and U66U144(tU66U144Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U66U145(tU66U145Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U66U146(tU66U146Out,~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U66U147(tU66U147Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U66U148(tU66U148Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:67====================
wire tU67U17Out;
wire tU67U123Out;
wire tU67U129Out;
wire tU67U13Out;
wire tU67U115Out;
wire tU67U120Out;
wire tU67U16Out;
wire tU67U12Out;
wire tU67U15Out;
wire tU67U19Out;
wire tU67U126Out;
wire tU67U10Out;
wire tU67U00Out;
wire tU67U128Out;
wire tU67U111Out;
wire tU67U11Out;
wire tU67U122Out;
wire tU67U121Out;
wire tU67U18Out;
wire tU67U112Out;
wire tU67U127Out;
wire tU67U116Out;
wire tU67U124Out;
wire tU67U113Out;
wire tU67U125Out;
wire tU67U119Out;
wire tU67U110Out;
wire tU67U118Out;
wire tU67U14Out;
wire tU67U114Out;
wire tU67U117Out;
or U67U00(tU67U00Out,tU67U10Out,tU67U11Out,tU67U12Out,tU67U13Out,tU67U14Out,tU67U15Out,tU67U16Out,tU67U17Out,tU67U18Out,tU67U19Out,tU67U110Out,tU67U111Out,tU67U112Out,tU67U113Out,tU67U114Out,tU67U115Out,tU67U116Out,tU67U117Out,tU67U118Out,tU67U119Out,tU67U120Out,tU67U121Out,tU67U122Out,tU67U123Out,tU67U124Out,tU67U125Out,tU67U126Out,tU67U127Out,tU67U128Out,tU67U129Out);
and U67U10(tU67U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U67U11(tU67U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U67U12(tU67U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U67U13(tU67U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U67U14(tU67U14Out,counter[1],~counter[2],counter[4],counter[5]);
and U67U15(tU67U15Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U67U16(tU67U16Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U67U17(tU67U17Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U67U18(tU67U18Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U67U19(tU67U19Out,~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U67U110(tU67U110Out,~counter[1],~counter[3],counter[4],counter[5]);
and U67U111(tU67U111Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U67U112(tU67U112Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U67U113(tU67U113Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U67U114(tU67U114Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U67U115(tU67U115Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U67U116(tU67U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U67U117(tU67U117Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U67U118(tU67U118Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U67U119(tU67U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U67U120(tU67U120Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U67U121(tU67U121Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U67U122(tU67U122Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U67U123(tU67U123Out,~counter[0],counter[2],counter[3],counter[5]);
and U67U124(tU67U124Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U67U125(tU67U125Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U67U126(tU67U126Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U67U127(tU67U127Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U67U128(tU67U128Out,~counter[1],counter[2],counter[3],counter[5]);
and U67U129(tU67U129Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:68====================
wire tU68U14Out;
wire tU68U122Out;
wire tU68U117Out;
wire tU68U10Out;
wire tU68U121Out;
wire tU68U114Out;
wire tU68U13Out;
wire tU68U18Out;
wire tU68U19Out;
wire tU68U129Out;
wire tU68U126Out;
wire tU68U16Out;
wire tU68U119Out;
wire tU68U112Out;
wire tU68U113Out;
wire tU68U110Out;
wire tU68U118Out;
wire tU68U00Out;
wire tU68U128Out;
wire tU68U127Out;
wire tU68U124Out;
wire tU68U111Out;
wire tU68U11Out;
wire tU68U116Out;
wire tU68U120Out;
wire tU68U123Out;
wire tU68U17Out;
wire tU68U12Out;
wire tU68U115Out;
wire tU68U15Out;
wire tU68U125Out;
or U68U00(tU68U00Out,tU68U10Out,tU68U11Out,tU68U12Out,tU68U13Out,tU68U14Out,tU68U15Out,tU68U16Out,tU68U17Out,tU68U18Out,tU68U19Out,tU68U110Out,tU68U111Out,tU68U112Out,tU68U113Out,tU68U114Out,tU68U115Out,tU68U116Out,tU68U117Out,tU68U118Out,tU68U119Out,tU68U120Out,tU68U121Out,tU68U122Out,tU68U123Out,tU68U124Out,tU68U125Out,tU68U126Out,tU68U127Out,tU68U128Out,tU68U129Out);
and U68U10(tU68U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U68U11(tU68U11Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U68U12(tU68U12Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U68U13(tU68U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U68U14(tU68U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U68U15(tU68U15Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U68U16(tU68U16Out,~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U68U17(tU68U17Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U68U18(tU68U18Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U68U19(tU68U19Out,~counter[1],~counter[3],counter[4],counter[5]);
and U68U110(tU68U110Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U68U111(tU68U111Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U68U112(tU68U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U68U113(tU68U113Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U68U114(tU68U114Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U68U115(tU68U115Out,~counter[0],~counter[1],~counter[3],~counter[4],~counter[5],counter[6]);
and U68U116(tU68U116Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U68U117(tU68U117Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U68U118(tU68U118Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U68U119(tU68U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U68U120(tU68U120Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U68U121(tU68U121Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U68U122(tU68U122Out,~counter[0],counter[2],counter[3],counter[5]);
and U68U123(tU68U123Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U68U124(tU68U124Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U68U125(tU68U125Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U68U126(tU68U126Out,~counter[1],counter[2],counter[3],counter[5]);
and U68U127(tU68U127Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U68U128(tU68U128Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U68U129(tU68U129Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:69====================
wire tU69U120Out;
wire tU69U114Out;
wire tU69U17Out;
wire tU69U118Out;
wire tU69U110Out;
wire tU69U115Out;
wire tU69U117Out;
wire tU69U111Out;
wire tU69U19Out;
wire tU69U10Out;
wire tU69U116Out;
wire tU69U121Out;
wire tU69U00Out;
wire tU69U123Out;
wire tU69U16Out;
wire tU69U13Out;
wire tU69U12Out;
wire tU69U113Out;
wire tU69U15Out;
wire tU69U122Out;
wire tU69U112Out;
wire tU69U119Out;
wire tU69U11Out;
wire tU69U18Out;
wire tU69U14Out;
or U69U00(tU69U00Out,tU69U10Out,tU69U11Out,tU69U12Out,tU69U13Out,tU69U14Out,tU69U15Out,tU69U16Out,tU69U17Out,tU69U18Out,tU69U19Out,tU69U110Out,tU69U111Out,tU69U112Out,tU69U113Out,tU69U114Out,tU69U115Out,tU69U116Out,tU69U117Out,tU69U118Out,tU69U119Out,tU69U120Out,tU69U121Out,tU69U122Out,tU69U123Out);
and U69U10(tU69U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U69U11(tU69U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U69U12(tU69U12Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U69U13(tU69U13Out,~counter[1],~counter[3],~counter[4],~counter[5],counter[6]);
and U69U14(tU69U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U69U15(tU69U15Out,counter[1],~counter[2],counter[4],counter[5]);
and U69U16(tU69U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U69U17(tU69U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U69U18(tU69U18Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U69U19(tU69U19Out,~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U69U110(tU69U110Out,~counter[1],~counter[3],counter[4],counter[5]);
and U69U111(tU69U111Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U69U112(tU69U112Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U69U113(tU69U113Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U69U114(tU69U114Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U69U115(tU69U115Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U69U116(tU69U116Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U69U117(tU69U117Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U69U118(tU69U118Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U69U119(tU69U119Out,~counter[0],counter[2],counter[3],counter[5]);
and U69U120(tU69U120Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U69U121(tU69U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U69U122(tU69U122Out,~counter[1],counter[2],counter[3],counter[5]);
and U69U123(tU69U123Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:70====================
wire tU70U19Out;
wire tU70U118Out;
wire tU70U11Out;
wire tU70U132Out;
wire tU70U125Out;
wire tU70U123Out;
wire tU70U140Out;
wire tU70U122Out;
wire tU70U13Out;
wire tU70U121Out;
wire tU70U131Out;
wire tU70U144Out;
wire tU70U147Out;
wire tU70U14Out;
wire tU70U137Out;
wire tU70U148Out;
wire tU70U135Out;
wire tU70U145Out;
wire tU70U146Out;
wire tU70U00Out;
wire tU70U12Out;
wire tU70U120Out;
wire tU70U136Out;
wire tU70U141Out;
wire tU70U114Out;
wire tU70U128Out;
wire tU70U119Out;
wire tU70U129Out;
wire tU70U116Out;
wire tU70U115Out;
wire tU70U139Out;
wire tU70U18Out;
wire tU70U17Out;
wire tU70U117Out;
wire tU70U127Out;
wire tU70U110Out;
wire tU70U134Out;
wire tU70U138Out;
wire tU70U149Out;
wire tU70U126Out;
wire tU70U143Out;
wire tU70U124Out;
wire tU70U112Out;
wire tU70U15Out;
wire tU70U113Out;
wire tU70U130Out;
wire tU70U133Out;
wire tU70U16Out;
wire tU70U142Out;
wire tU70U10Out;
wire tU70U111Out;
or U70U00(tU70U00Out,tU70U10Out,tU70U11Out,tU70U12Out,tU70U13Out,tU70U14Out,tU70U15Out,tU70U16Out,tU70U17Out,tU70U18Out,tU70U19Out,tU70U110Out,tU70U111Out,tU70U112Out,tU70U113Out,tU70U114Out,tU70U115Out,tU70U116Out,tU70U117Out,tU70U118Out,tU70U119Out,tU70U120Out,tU70U121Out,tU70U122Out,tU70U123Out,tU70U124Out,tU70U125Out,tU70U126Out,tU70U127Out,tU70U128Out,tU70U129Out,tU70U130Out,tU70U131Out,tU70U132Out,tU70U133Out,tU70U134Out,tU70U135Out,tU70U136Out,tU70U137Out,tU70U138Out,tU70U139Out,tU70U140Out,tU70U141Out,tU70U142Out,tU70U143Out,tU70U144Out,tU70U145Out,tU70U146Out,tU70U147Out,tU70U148Out,tU70U149Out);
and U70U10(tU70U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U70U11(tU70U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U70U12(tU70U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U70U13(tU70U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U70U14(tU70U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U70U15(tU70U15Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U70U16(tU70U16Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U70U17(tU70U17Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U70U18(tU70U18Out,~counter[1],~counter[3],~counter[4],~counter[5],counter[6]);
and U70U19(tU70U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U70U110(tU70U110Out,counter[1],~counter[2],counter[4],counter[5]);
and U70U111(tU70U111Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U70U112(tU70U112Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U70U113(tU70U113Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U70U114(tU70U114Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U70U115(tU70U115Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U70U116(tU70U116Out,~counter[2],~counter[3],~counter[4],~counter[5],counter[6]);
and U70U117(tU70U117Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U70U118(tU70U118Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U70U119(tU70U119Out,~counter[1],~counter[3],counter[4],counter[5]);
and U70U120(tU70U120Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U70U121(tU70U121Out,~counter[0],~counter[3],~counter[4],~counter[5],counter[6]);
and U70U122(tU70U122Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U70U123(tU70U123Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U70U124(tU70U124Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U70U125(tU70U125Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U70U126(tU70U126Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U70U127(tU70U127Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U70U128(tU70U128Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U70U129(tU70U129Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U70U130(tU70U130Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U70U131(tU70U131Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U70U132(tU70U132Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U70U133(tU70U133Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U70U134(tU70U134Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U70U135(tU70U135Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U70U136(tU70U136Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U70U137(tU70U137Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U70U138(tU70U138Out,~counter[0],counter[2],counter[3],counter[5]);
and U70U139(tU70U139Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U70U140(tU70U140Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U70U141(tU70U141Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U70U142(tU70U142Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U70U143(tU70U143Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U70U144(tU70U144Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U70U145(tU70U145Out,~counter[1],counter[2],counter[3],counter[5]);
and U70U146(tU70U146Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U70U147(tU70U147Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U70U148(tU70U148Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U70U149(tU70U149Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:71====================
wire tU71U14Out;
wire tU71U126Out;
wire tU71U00Out;
wire tU71U13Out;
wire tU71U119Out;
wire tU71U11Out;
wire tU71U17Out;
wire tU71U118Out;
wire tU71U127Out;
wire tU71U18Out;
wire tU71U15Out;
wire tU71U117Out;
wire tU71U120Out;
wire tU71U125Out;
wire tU71U116Out;
wire tU71U123Out;
wire tU71U16Out;
wire tU71U12Out;
wire tU71U113Out;
wire tU71U121Out;
wire tU71U122Out;
wire tU71U114Out;
wire tU71U124Out;
wire tU71U115Out;
wire tU71U10Out;
wire tU71U111Out;
wire tU71U110Out;
wire tU71U19Out;
wire tU71U112Out;
or U71U00(tU71U00Out,tU71U10Out,tU71U11Out,tU71U12Out,tU71U13Out,tU71U14Out,tU71U15Out,tU71U16Out,tU71U17Out,tU71U18Out,tU71U19Out,tU71U110Out,tU71U111Out,tU71U112Out,tU71U113Out,tU71U114Out,tU71U115Out,tU71U116Out,tU71U117Out,tU71U118Out,tU71U119Out,tU71U120Out,tU71U121Out,tU71U122Out,tU71U123Out,tU71U124Out,tU71U125Out,tU71U126Out,tU71U127Out);
and U71U10(tU71U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U71U11(tU71U11Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U71U12(tU71U12Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U71U13(tU71U13Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U71U14(tU71U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U71U15(tU71U15Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U71U16(tU71U16Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U71U17(tU71U17Out,counter[1],~counter[2],counter[4],counter[5]);
and U71U18(tU71U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U71U19(tU71U19Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U71U110(tU71U110Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U71U111(tU71U111Out,~counter[1],~counter[3],counter[4],counter[5]);
and U71U112(tU71U112Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U71U113(tU71U113Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U71U114(tU71U114Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U71U115(tU71U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U71U116(tU71U116Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U71U117(tU71U117Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U71U118(tU71U118Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U71U119(tU71U119Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U71U120(tU71U120Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U71U121(tU71U121Out,~counter[0],counter[2],counter[3],counter[5]);
and U71U122(tU71U122Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U71U123(tU71U123Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U71U124(tU71U124Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U71U125(tU71U125Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U71U126(tU71U126Out,~counter[1],counter[2],counter[3],counter[5]);
and U71U127(tU71U127Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:72====================
wire tU72U146Out;
wire tU72U13Out;
wire tU72U142Out;
wire tU72U10Out;
wire tU72U112Out;
wire tU72U115Out;
wire tU72U114Out;
wire tU72U117Out;
wire tU72U132Out;
wire tU72U133Out;
wire tU72U110Out;
wire tU72U122Out;
wire tU72U19Out;
wire tU72U11Out;
wire tU72U135Out;
wire tU72U139Out;
wire tU72U119Out;
wire tU72U121Out;
wire tU72U130Out;
wire tU72U143Out;
wire tU72U137Out;
wire tU72U123Out;
wire tU72U126Out;
wire tU72U120Out;
wire tU72U12Out;
wire tU72U128Out;
wire tU72U148Out;
wire tU72U147Out;
wire tU72U136Out;
wire tU72U125Out;
wire tU72U18Out;
wire tU72U116Out;
wire tU72U113Out;
wire tU72U17Out;
wire tU72U129Out;
wire tU72U138Out;
wire tU72U141Out;
wire tU72U145Out;
wire tU72U140Out;
wire tU72U127Out;
wire tU72U131Out;
wire tU72U144Out;
wire tU72U16Out;
wire tU72U118Out;
wire tU72U14Out;
wire tU72U00Out;
wire tU72U124Out;
wire tU72U111Out;
wire tU72U15Out;
wire tU72U134Out;
or U72U00(tU72U00Out,tU72U10Out,tU72U11Out,tU72U12Out,tU72U13Out,tU72U14Out,tU72U15Out,tU72U16Out,tU72U17Out,tU72U18Out,tU72U19Out,tU72U110Out,tU72U111Out,tU72U112Out,tU72U113Out,tU72U114Out,tU72U115Out,tU72U116Out,tU72U117Out,tU72U118Out,tU72U119Out,tU72U120Out,tU72U121Out,tU72U122Out,tU72U123Out,tU72U124Out,tU72U125Out,tU72U126Out,tU72U127Out,tU72U128Out,tU72U129Out,tU72U130Out,tU72U131Out,tU72U132Out,tU72U133Out,tU72U134Out,tU72U135Out,tU72U136Out,tU72U137Out,tU72U138Out,tU72U139Out,tU72U140Out,tU72U141Out,tU72U142Out,tU72U143Out,tU72U144Out,tU72U145Out,tU72U146Out,tU72U147Out,tU72U148Out);
and U72U10(tU72U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U72U11(tU72U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U72U12(tU72U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U72U13(tU72U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U72U14(tU72U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U72U15(tU72U15Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U72U16(tU72U16Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U72U17(tU72U17Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U72U18(tU72U18Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U72U19(tU72U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U72U110(tU72U110Out,counter[1],~counter[2],counter[4],counter[5]);
and U72U111(tU72U111Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U72U112(tU72U112Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U72U113(tU72U113Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U72U114(tU72U114Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U72U115(tU72U115Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U72U116(tU72U116Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U72U117(tU72U117Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U72U118(tU72U118Out,~counter[1],~counter[3],counter[4],counter[5]);
and U72U119(tU72U119Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U72U120(tU72U120Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U72U121(tU72U121Out,~counter[0],~counter[1],~counter[2],~counter[4],~counter[5],counter[6]);
and U72U122(tU72U122Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U72U123(tU72U123Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U72U124(tU72U124Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U72U125(tU72U125Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U72U126(tU72U126Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U72U127(tU72U127Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U72U128(tU72U128Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U72U129(tU72U129Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U72U130(tU72U130Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U72U131(tU72U131Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U72U132(tU72U132Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U72U133(tU72U133Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U72U134(tU72U134Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U72U135(tU72U135Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U72U136(tU72U136Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U72U137(tU72U137Out,~counter[0],counter[2],counter[3],counter[5]);
and U72U138(tU72U138Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U72U139(tU72U139Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U72U140(tU72U140Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U72U141(tU72U141Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U72U142(tU72U142Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U72U143(tU72U143Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U72U144(tU72U144Out,~counter[1],counter[2],counter[3],counter[5]);
and U72U145(tU72U145Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U72U146(tU72U146Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U72U147(tU72U147Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U72U148(tU72U148Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:73====================
wire tU73U111Out;
wire tU73U14Out;
wire tU73U13Out;
wire tU73U10Out;
wire tU73U110Out;
wire tU73U112Out;
wire tU73U18Out;
wire tU73U00Out;
wire tU73U113Out;
wire tU73U116Out;
wire tU73U17Out;
wire tU73U16Out;
wire tU73U114Out;
wire tU73U15Out;
wire tU73U19Out;
wire tU73U11Out;
wire tU73U115Out;
wire tU73U12Out;
or U73U00(tU73U00Out,tU73U10Out,tU73U11Out,tU73U12Out,tU73U13Out,tU73U14Out,tU73U15Out,tU73U16Out,tU73U17Out,tU73U18Out,tU73U19Out,tU73U110Out,tU73U111Out,tU73U112Out,tU73U113Out,tU73U114Out,tU73U115Out,tU73U116Out);
and U73U10(tU73U10Out,~counter[1],~counter[2],~counter[4],~counter[5],counter[6]);
and U73U11(tU73U11Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U73U12(tU73U12Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U73U13(tU73U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U73U14(tU73U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U73U15(tU73U15Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U73U16(tU73U16Out,~counter[1],~counter[3],counter[4],counter[5]);
and U73U17(tU73U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U73U18(tU73U18Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U73U19(tU73U19Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U73U110(tU73U110Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U73U111(tU73U111Out,~counter[0],counter[2],counter[3],counter[5]);
and U73U112(tU73U112Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U73U113(tU73U113Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U73U114(tU73U114Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U73U115(tU73U115Out,~counter[1],counter[2],counter[3],counter[5]);
and U73U116(tU73U116Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:74====================
wire tU74U122Out;
wire tU74U128Out;
wire tU74U123Out;
wire tU74U12Out;
wire tU74U10Out;
wire tU74U00Out;
wire tU74U118Out;
wire tU74U11Out;
wire tU74U112Out;
wire tU74U115Out;
wire tU74U126Out;
wire tU74U15Out;
wire tU74U17Out;
wire tU74U119Out;
wire tU74U129Out;
wire tU74U120Out;
wire tU74U14Out;
wire tU74U125Out;
wire tU74U132Out;
wire tU74U133Out;
wire tU74U121Out;
wire tU74U16Out;
wire tU74U131Out;
wire tU74U117Out;
wire tU74U124Out;
wire tU74U19Out;
wire tU74U127Out;
wire tU74U18Out;
wire tU74U130Out;
wire tU74U113Out;
wire tU74U114Out;
wire tU74U111Out;
wire tU74U116Out;
wire tU74U13Out;
wire tU74U110Out;
wire tU74U134Out;
or U74U00(tU74U00Out,tU74U10Out,tU74U11Out,tU74U12Out,tU74U13Out,tU74U14Out,tU74U15Out,tU74U16Out,tU74U17Out,tU74U18Out,tU74U19Out,tU74U110Out,tU74U111Out,tU74U112Out,tU74U113Out,tU74U114Out,tU74U115Out,tU74U116Out,tU74U117Out,tU74U118Out,tU74U119Out,tU74U120Out,tU74U121Out,tU74U122Out,tU74U123Out,tU74U124Out,tU74U125Out,tU74U126Out,tU74U127Out,tU74U128Out,tU74U129Out,tU74U130Out,tU74U131Out,tU74U132Out,tU74U133Out,tU74U134Out);
and U74U10(tU74U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U74U11(tU74U11Out,~counter[1],~counter[2],~counter[4],~counter[5],counter[6]);
and U74U12(tU74U12Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U74U13(tU74U13Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U74U14(tU74U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U74U15(tU74U15Out,counter[1],~counter[2],counter[4],counter[5]);
and U74U16(tU74U16Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U74U17(tU74U17Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U74U18(tU74U18Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U74U19(tU74U19Out,counter[0],counter[3],counter[4],~counter[5],~counter[6]);
and U74U110(tU74U110Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U74U111(tU74U111Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U74U112(tU74U112Out,~counter[1],~counter[3],counter[4],counter[5]);
and U74U113(tU74U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U74U114(tU74U114Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U74U115(tU74U115Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U74U116(tU74U116Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U74U117(tU74U117Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U74U118(tU74U118Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U74U119(tU74U119Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U74U120(tU74U120Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U74U121(tU74U121Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U74U122(tU74U122Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U74U123(tU74U123Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U74U124(tU74U124Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U74U125(tU74U125Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U74U126(tU74U126Out,~counter[0],counter[2],counter[3],counter[5]);
and U74U127(tU74U127Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U74U128(tU74U128Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U74U129(tU74U129Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U74U130(tU74U130Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U74U131(tU74U131Out,~counter[1],counter[2],counter[3],counter[5]);
and U74U132(tU74U132Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U74U133(tU74U133Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U74U134(tU74U134Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:75====================
wire tU75U12Out;
wire tU75U123Out;
wire tU75U121Out;
wire tU75U126Out;
wire tU75U119Out;
wire tU75U18Out;
wire tU75U127Out;
wire tU75U110Out;
wire tU75U125Out;
wire tU75U115Out;
wire tU75U16Out;
wire tU75U118Out;
wire tU75U122Out;
wire tU75U128Out;
wire tU75U13Out;
wire tU75U112Out;
wire tU75U11Out;
wire tU75U116Out;
wire tU75U111Out;
wire tU75U113Out;
wire tU75U120Out;
wire tU75U17Out;
wire tU75U117Out;
wire tU75U10Out;
wire tU75U124Out;
wire tU75U14Out;
wire tU75U00Out;
wire tU75U19Out;
wire tU75U15Out;
wire tU75U114Out;
or U75U00(tU75U00Out,tU75U10Out,tU75U11Out,tU75U12Out,tU75U13Out,tU75U14Out,tU75U15Out,tU75U16Out,tU75U17Out,tU75U18Out,tU75U19Out,tU75U110Out,tU75U111Out,tU75U112Out,tU75U113Out,tU75U114Out,tU75U115Out,tU75U116Out,tU75U117Out,tU75U118Out,tU75U119Out,tU75U120Out,tU75U121Out,tU75U122Out,tU75U123Out,tU75U124Out,tU75U125Out,tU75U126Out,tU75U127Out,tU75U128Out);
and U75U10(tU75U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U75U11(tU75U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U75U12(tU75U12Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U75U13(tU75U13Out,~counter[2],~counter[4],~counter[5],counter[6]);
and U75U14(tU75U14Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U75U15(tU75U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U75U16(tU75U16Out,counter[1],~counter[2],counter[4],counter[5]);
and U75U17(tU75U17Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U75U18(tU75U18Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U75U19(tU75U19Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U75U110(tU75U110Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U75U111(tU75U111Out,~counter[1],~counter[3],counter[4],counter[5]);
and U75U112(tU75U112Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U75U113(tU75U113Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U75U114(tU75U114Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U75U115(tU75U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U75U116(tU75U116Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U75U117(tU75U117Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U75U118(tU75U118Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U75U119(tU75U119Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U75U120(tU75U120Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U75U121(tU75U121Out,~counter[0],counter[2],counter[3],counter[5]);
and U75U122(tU75U122Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U75U123(tU75U123Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U75U124(tU75U124Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U75U125(tU75U125Out,~counter[1],counter[2],counter[3],counter[5]);
and U75U126(tU75U126Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U75U127(tU75U127Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U75U128(tU75U128Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:76====================
wire tU76U129Out;
wire tU76U140Out;
wire tU76U126Out;
wire tU76U125Out;
wire tU76U143Out;
wire tU76U18Out;
wire tU76U14Out;
wire tU76U127Out;
wire tU76U00Out;
wire tU76U12Out;
wire tU76U114Out;
wire tU76U112Out;
wire tU76U119Out;
wire tU76U128Out;
wire tU76U139Out;
wire tU76U115Out;
wire tU76U130Out;
wire tU76U17Out;
wire tU76U145Out;
wire tU76U116Out;
wire tU76U141Out;
wire tU76U122Out;
wire tU76U136Out;
wire tU76U16Out;
wire tU76U144Out;
wire tU76U19Out;
wire tU76U124Out;
wire tU76U131Out;
wire tU76U134Out;
wire tU76U146Out;
wire tU76U135Out;
wire tU76U111Out;
wire tU76U13Out;
wire tU76U120Out;
wire tU76U138Out;
wire tU76U10Out;
wire tU76U118Out;
wire tU76U137Out;
wire tU76U110Out;
wire tU76U132Out;
wire tU76U15Out;
wire tU76U113Out;
wire tU76U123Out;
wire tU76U121Out;
wire tU76U142Out;
wire tU76U117Out;
wire tU76U133Out;
wire tU76U11Out;
or U76U00(tU76U00Out,tU76U10Out,tU76U11Out,tU76U12Out,tU76U13Out,tU76U14Out,tU76U15Out,tU76U16Out,tU76U17Out,tU76U18Out,tU76U19Out,tU76U110Out,tU76U111Out,tU76U112Out,tU76U113Out,tU76U114Out,tU76U115Out,tU76U116Out,tU76U117Out,tU76U118Out,tU76U119Out,tU76U120Out,tU76U121Out,tU76U122Out,tU76U123Out,tU76U124Out,tU76U125Out,tU76U126Out,tU76U127Out,tU76U128Out,tU76U129Out,tU76U130Out,tU76U131Out,tU76U132Out,tU76U133Out,tU76U134Out,tU76U135Out,tU76U136Out,tU76U137Out,tU76U138Out,tU76U139Out,tU76U140Out,tU76U141Out,tU76U142Out,tU76U143Out,tU76U144Out,tU76U145Out,tU76U146Out);
and U76U10(tU76U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U76U11(tU76U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U76U12(tU76U12Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U76U13(tU76U13Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U76U14(tU76U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U76U15(tU76U15Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U76U16(tU76U16Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U76U17(tU76U17Out,~counter[2],~counter[4],~counter[5],counter[6]);
and U76U18(tU76U18Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U76U19(tU76U19Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U76U110(tU76U110Out,~counter[0],~counter[1],~counter[4],~counter[5],counter[6]);
and U76U111(tU76U111Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U76U112(tU76U112Out,counter[1],~counter[2],counter[4],counter[5]);
and U76U113(tU76U113Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U76U114(tU76U114Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U76U115(tU76U115Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U76U116(tU76U116Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U76U117(tU76U117Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U76U118(tU76U118Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U76U119(tU76U119Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U76U120(tU76U120Out,~counter[1],~counter[3],counter[4],counter[5]);
and U76U121(tU76U121Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U76U122(tU76U122Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U76U123(tU76U123Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U76U124(tU76U124Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U76U125(tU76U125Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U76U126(tU76U126Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U76U127(tU76U127Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U76U128(tU76U128Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U76U129(tU76U129Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U76U130(tU76U130Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U76U131(tU76U131Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U76U132(tU76U132Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U76U133(tU76U133Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U76U134(tU76U134Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U76U135(tU76U135Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U76U136(tU76U136Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U76U137(tU76U137Out,~counter[0],counter[2],counter[3],counter[5]);
and U76U138(tU76U138Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U76U139(tU76U139Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U76U140(tU76U140Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U76U141(tU76U141Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U76U142(tU76U142Out,~counter[1],counter[2],counter[3],counter[5]);
and U76U143(tU76U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U76U144(tU76U144Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U76U145(tU76U145Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U76U146(tU76U146Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:77====================
wire tU77U13Out;
wire tU77U113Out;
wire tU77U117Out;
wire tU77U19Out;
wire tU77U121Out;
wire tU77U125Out;
wire tU77U124Out;
wire tU77U110Out;
wire tU77U10Out;
wire tU77U12Out;
wire tU77U119Out;
wire tU77U116Out;
wire tU77U114Out;
wire tU77U126Out;
wire tU77U127Out;
wire tU77U15Out;
wire tU77U11Out;
wire tU77U17Out;
wire tU77U112Out;
wire tU77U118Out;
wire tU77U115Out;
wire tU77U16Out;
wire tU77U111Out;
wire tU77U18Out;
wire tU77U123Out;
wire tU77U14Out;
wire tU77U122Out;
wire tU77U120Out;
wire tU77U128Out;
wire tU77U00Out;
or U77U00(tU77U00Out,tU77U10Out,tU77U11Out,tU77U12Out,tU77U13Out,tU77U14Out,tU77U15Out,tU77U16Out,tU77U17Out,tU77U18Out,tU77U19Out,tU77U110Out,tU77U111Out,tU77U112Out,tU77U113Out,tU77U114Out,tU77U115Out,tU77U116Out,tU77U117Out,tU77U118Out,tU77U119Out,tU77U120Out,tU77U121Out,tU77U122Out,tU77U123Out,tU77U124Out,tU77U125Out,tU77U126Out,tU77U127Out,tU77U128Out);
and U77U10(tU77U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U77U11(tU77U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U77U12(tU77U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U77U13(tU77U13Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U77U14(tU77U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U77U15(tU77U15Out,~counter[2],~counter[4],~counter[5],counter[6]);
and U77U16(tU77U16Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U77U17(tU77U17Out,~counter[0],~counter[1],~counter[4],~counter[5],counter[6]);
and U77U18(tU77U18Out,counter[1],~counter[2],counter[4],counter[5]);
and U77U19(tU77U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U77U110(tU77U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U77U111(tU77U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U77U112(tU77U112Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U77U113(tU77U113Out,~counter[1],~counter[3],counter[4],counter[5]);
and U77U114(tU77U114Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U77U115(tU77U115Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U77U116(tU77U116Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U77U117(tU77U117Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U77U118(tU77U118Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U77U119(tU77U119Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U77U120(tU77U120Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U77U121(tU77U121Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U77U122(tU77U122Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U77U123(tU77U123Out,~counter[0],counter[2],counter[3],counter[5]);
and U77U124(tU77U124Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U77U125(tU77U125Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U77U126(tU77U126Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U77U127(tU77U127Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U77U128(tU77U128Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:78====================
wire tU78U146Out;
wire tU78U114Out;
wire tU78U12Out;
wire tU78U143Out;
wire tU78U11Out;
wire tU78U10Out;
wire tU78U132Out;
wire tU78U129Out;
wire tU78U119Out;
wire tU78U138Out;
wire tU78U121Out;
wire tU78U127Out;
wire tU78U140Out;
wire tU78U128Out;
wire tU78U136Out;
wire tU78U118Out;
wire tU78U115Out;
wire tU78U123Out;
wire tU78U17Out;
wire tU78U14Out;
wire tU78U137Out;
wire tU78U00Out;
wire tU78U112Out;
wire tU78U111Out;
wire tU78U134Out;
wire tU78U135Out;
wire tU78U117Out;
wire tU78U126Out;
wire tU78U130Out;
wire tU78U141Out;
wire tU78U15Out;
wire tU78U18Out;
wire tU78U110Out;
wire tU78U125Out;
wire tU78U120Out;
wire tU78U144Out;
wire tU78U113Out;
wire tU78U131Out;
wire tU78U13Out;
wire tU78U16Out;
wire tU78U145Out;
wire tU78U142Out;
wire tU78U124Out;
wire tU78U139Out;
wire tU78U19Out;
wire tU78U116Out;
wire tU78U133Out;
wire tU78U122Out;
or U78U00(tU78U00Out,tU78U10Out,tU78U11Out,tU78U12Out,tU78U13Out,tU78U14Out,tU78U15Out,tU78U16Out,tU78U17Out,tU78U18Out,tU78U19Out,tU78U110Out,tU78U111Out,tU78U112Out,tU78U113Out,tU78U114Out,tU78U115Out,tU78U116Out,tU78U117Out,tU78U118Out,tU78U119Out,tU78U120Out,tU78U121Out,tU78U122Out,tU78U123Out,tU78U124Out,tU78U125Out,tU78U126Out,tU78U127Out,tU78U128Out,tU78U129Out,tU78U130Out,tU78U131Out,tU78U132Out,tU78U133Out,tU78U134Out,tU78U135Out,tU78U136Out,tU78U137Out,tU78U138Out,tU78U139Out,tU78U140Out,tU78U141Out,tU78U142Out,tU78U143Out,tU78U144Out,tU78U145Out,tU78U146Out);
and U78U10(tU78U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U78U11(tU78U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U78U12(tU78U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U78U13(tU78U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U78U14(tU78U14Out,~counter[3],~counter[4],~counter[5],counter[6]);
and U78U15(tU78U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U78U16(tU78U16Out,~counter[2],~counter[4],~counter[5],counter[6]);
and U78U17(tU78U17Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U78U18(tU78U18Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U78U19(tU78U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U78U110(tU78U110Out,counter[1],~counter[2],counter[4],counter[5]);
and U78U111(tU78U111Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U78U112(tU78U112Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U78U113(tU78U113Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U78U114(tU78U114Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U78U115(tU78U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U78U116(tU78U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U78U117(tU78U117Out,~counter[1],~counter[3],counter[4],counter[5]);
and U78U118(tU78U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U78U119(tU78U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U78U120(tU78U120Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U78U121(tU78U121Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U78U122(tU78U122Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U78U123(tU78U123Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U78U124(tU78U124Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U78U125(tU78U125Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U78U126(tU78U126Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U78U127(tU78U127Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U78U128(tU78U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U78U129(tU78U129Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U78U130(tU78U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U78U131(tU78U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U78U132(tU78U132Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U78U133(tU78U133Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U78U134(tU78U134Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U78U135(tU78U135Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U78U136(tU78U136Out,~counter[0],counter[2],counter[3],counter[5]);
and U78U137(tU78U137Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U78U138(tU78U138Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U78U139(tU78U139Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U78U140(tU78U140Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U78U141(tU78U141Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U78U142(tU78U142Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U78U143(tU78U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U78U144(tU78U144Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U78U145(tU78U145Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U78U146(tU78U146Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:79====================
wire tU79U16Out;
wire tU79U13Out;
wire tU79U14Out;
wire tU79U112Out;
wire tU79U117Out;
wire tU79U115Out;
wire tU79U116Out;
wire tU79U10Out;
wire tU79U114Out;
wire tU79U00Out;
wire tU79U15Out;
wire tU79U11Out;
wire tU79U113Out;
wire tU79U12Out;
wire tU79U17Out;
wire tU79U111Out;
wire tU79U19Out;
wire tU79U18Out;
wire tU79U110Out;
or U79U00(tU79U00Out,tU79U10Out,tU79U11Out,tU79U12Out,tU79U13Out,tU79U14Out,tU79U15Out,tU79U16Out,tU79U17Out,tU79U18Out,tU79U19Out,tU79U110Out,tU79U111Out,tU79U112Out,tU79U113Out,tU79U114Out,tU79U115Out,tU79U116Out,tU79U117Out);
and U79U10(tU79U10Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U79U11(tU79U11Out,counter[1],~counter[2],counter[4],counter[5]);
and U79U12(tU79U12Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U79U13(tU79U13Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U79U14(tU79U14Out,~counter[1],~counter[3],counter[4],counter[5]);
and U79U15(tU79U15Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U79U16(tU79U16Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U79U17(tU79U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U79U18(tU79U18Out,~counter[4],~counter[5],counter[6]);
and U79U19(tU79U19Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U79U110(tU79U110Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U79U111(tU79U111Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U79U112(tU79U112Out,~counter[0],counter[2],counter[3],counter[5]);
and U79U113(tU79U113Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U79U114(tU79U114Out,~counter[0],~counter[1],~counter[2],counter[3],~counter[4],~counter[6]);
and U79U115(tU79U115Out,~counter[1],counter[2],counter[3],counter[5]);
and U79U116(tU79U116Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U79U117(tU79U117Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:80====================
wire tU80U119Out;
wire tU80U118Out;
wire tU80U17Out;
wire tU80U16Out;
wire tU80U120Out;
wire tU80U18Out;
wire tU80U122Out;
wire tU80U12Out;
wire tU80U15Out;
wire tU80U113Out;
wire tU80U121Out;
wire tU80U13Out;
wire tU80U19Out;
wire tU80U114Out;
wire tU80U115Out;
wire tU80U112Out;
wire tU80U116Out;
wire tU80U111Out;
wire tU80U10Out;
wire tU80U00Out;
wire tU80U117Out;
wire tU80U110Out;
wire tU80U11Out;
wire tU80U14Out;
or U80U00(tU80U00Out,tU80U10Out,tU80U11Out,tU80U12Out,tU80U13Out,tU80U14Out,tU80U15Out,tU80U16Out,tU80U17Out,tU80U18Out,tU80U19Out,tU80U110Out,tU80U111Out,tU80U112Out,tU80U113Out,tU80U114Out,tU80U115Out,tU80U116Out,tU80U117Out,tU80U118Out,tU80U119Out,tU80U120Out,tU80U121Out,tU80U122Out);
and U80U10(tU80U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U11(tU80U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U80U12(tU80U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U80U13(tU80U13Out,counter[5],counter[6]);
and U80U14(tU80U14Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U80U15(tU80U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U16(tU80U16Out,counter[2],counter[4],counter[6]);
and U80U17(tU80U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U80U18(tU80U18Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U80U19(tU80U19Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U110(tU80U110Out,~counter[1],~counter[2],counter[3],counter[4],counter[6]);
and U80U111(tU80U111Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U112(tU80U112Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U80U113(tU80U113Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U114(tU80U114Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U80U115(tU80U115Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U116(tU80U116Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U80U117(tU80U117Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U80U118(tU80U118Out,counter[0],~counter[2],~counter[3],counter[4],counter[6]);
and U80U119(tU80U119Out,counter[1],~counter[2],counter[4],counter[6]);
and U80U120(tU80U120Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U80U121(tU80U121Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U80U122(tU80U122Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);

//====================Truthtable Variable:81====================
wire tU81U13Out;
wire tU81U110Out;
wire tU81U11Out;
wire tU81U19Out;
wire tU81U18Out;
wire tU81U111Out;
wire tU81U10Out;
wire tU81U12Out;
wire tU81U16Out;
wire tU81U17Out;
wire tU81U14Out;
wire tU81U00Out;
wire tU81U15Out;
wire tU81U112Out;
or U81U00(tU81U00Out,tU81U10Out,tU81U11Out,tU81U12Out,tU81U13Out,tU81U14Out,tU81U15Out,tU81U16Out,tU81U17Out,tU81U18Out,tU81U19Out,tU81U110Out,tU81U111Out,tU81U112Out);
and U81U10(tU81U10Out,counter[1],~counter[2],counter[4],counter[5]);
and U81U11(tU81U11Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U81U12(tU81U12Out,~counter[1],~counter[3],counter[4],counter[5]);
and U81U13(tU81U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U81U14(tU81U14Out,~counter[4],~counter[5],counter[6]);
and U81U15(tU81U15Out,~counter[1],~counter[2],~counter[3],~counter[5],counter[6]);
and U81U16(tU81U16Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U81U17(tU81U17Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U81U18(tU81U18Out,~counter[0],counter[2],counter[3],counter[5]);
and U81U19(tU81U19Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U81U110(tU81U110Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U81U111(tU81U111Out,~counter[1],counter[2],counter[3],counter[5]);
and U81U112(tU81U112Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:82====================
wire tU82U141Out;
wire tU82U17Out;
wire tU82U122Out;
wire tU82U138Out;
wire tU82U140Out;
wire tU82U112Out;
wire tU82U124Out;
wire tU82U128Out;
wire tU82U132Out;
wire tU82U16Out;
wire tU82U131Out;
wire tU82U130Out;
wire tU82U129Out;
wire tU82U136Out;
wire tU82U135Out;
wire tU82U139Out;
wire tU82U145Out;
wire tU82U12Out;
wire tU82U142Out;
wire tU82U118Out;
wire tU82U11Out;
wire tU82U00Out;
wire tU82U120Out;
wire tU82U111Out;
wire tU82U14Out;
wire tU82U110Out;
wire tU82U115Out;
wire tU82U15Out;
wire tU82U143Out;
wire tU82U117Out;
wire tU82U18Out;
wire tU82U126Out;
wire tU82U113Out;
wire tU82U19Out;
wire tU82U137Out;
wire tU82U123Out;
wire tU82U127Out;
wire tU82U119Out;
wire tU82U116Out;
wire tU82U10Out;
wire tU82U144Out;
wire tU82U134Out;
wire tU82U121Out;
wire tU82U13Out;
wire tU82U125Out;
wire tU82U133Out;
wire tU82U147Out;
wire tU82U146Out;
wire tU82U114Out;
or U82U00(tU82U00Out,tU82U10Out,tU82U11Out,tU82U12Out,tU82U13Out,tU82U14Out,tU82U15Out,tU82U16Out,tU82U17Out,tU82U18Out,tU82U19Out,tU82U110Out,tU82U111Out,tU82U112Out,tU82U113Out,tU82U114Out,tU82U115Out,tU82U116Out,tU82U117Out,tU82U118Out,tU82U119Out,tU82U120Out,tU82U121Out,tU82U122Out,tU82U123Out,tU82U124Out,tU82U125Out,tU82U126Out,tU82U127Out,tU82U128Out,tU82U129Out,tU82U130Out,tU82U131Out,tU82U132Out,tU82U133Out,tU82U134Out,tU82U135Out,tU82U136Out,tU82U137Out,tU82U138Out,tU82U139Out,tU82U140Out,tU82U141Out,tU82U142Out,tU82U143Out,tU82U144Out,tU82U145Out,tU82U146Out,tU82U147Out);
and U82U10(tU82U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U82U11(tU82U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U82U12(tU82U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U82U13(tU82U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U82U14(tU82U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U82U15(tU82U15Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U82U16(tU82U16Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U82U17(tU82U17Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U82U18(tU82U18Out,counter[1],~counter[2],counter[4],counter[5]);
and U82U19(tU82U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U82U110(tU82U110Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U82U111(tU82U111Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U82U112(tU82U112Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U82U113(tU82U113Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U82U114(tU82U114Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U82U115(tU82U115Out,~counter[1],~counter[3],counter[4],counter[5]);
and U82U116(tU82U116Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U82U117(tU82U117Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U82U118(tU82U118Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U82U119(tU82U119Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U82U120(tU82U120Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U82U121(tU82U121Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U82U122(tU82U122Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U82U123(tU82U123Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U82U124(tU82U124Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U82U125(tU82U125Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U82U126(tU82U126Out,~counter[4],~counter[5],counter[6]);
and U82U127(tU82U127Out,~counter[1],~counter[2],~counter[3],~counter[5],counter[6]);
and U82U128(tU82U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U82U129(tU82U129Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U82U130(tU82U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U82U131(tU82U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U82U132(tU82U132Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U82U133(tU82U133Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U82U134(tU82U134Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U82U135(tU82U135Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U82U136(tU82U136Out,~counter[0],~counter[2],~counter[3],~counter[5],counter[6]);
and U82U137(tU82U137Out,~counter[0],counter[2],counter[3],counter[5]);
and U82U138(tU82U138Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U82U139(tU82U139Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U82U140(tU82U140Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U82U141(tU82U141Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U82U142(tU82U142Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U82U143(tU82U143Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U82U144(tU82U144Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U82U145(tU82U145Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U82U146(tU82U146Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U82U147(tU82U147Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:83====================
wire tU83U15Out;
wire tU83U17Out;
wire tU83U19Out;
wire tU83U12Out;
wire tU83U115Out;
wire tU83U117Out;
wire tU83U119Out;
wire tU83U114Out;
wire tU83U11Out;
wire tU83U116Out;
wire tU83U10Out;
wire tU83U110Out;
wire tU83U113Out;
wire tU83U13Out;
wire tU83U00Out;
wire tU83U16Out;
wire tU83U120Out;
wire tU83U14Out;
wire tU83U118Out;
wire tU83U112Out;
wire tU83U111Out;
wire tU83U18Out;
or U83U00(tU83U00Out,tU83U10Out,tU83U11Out,tU83U12Out,tU83U13Out,tU83U14Out,tU83U15Out,tU83U16Out,tU83U17Out,tU83U18Out,tU83U19Out,tU83U110Out,tU83U111Out,tU83U112Out,tU83U113Out,tU83U114Out,tU83U115Out,tU83U116Out,tU83U117Out,tU83U118Out,tU83U119Out,tU83U120Out);
and U83U10(tU83U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U83U11(tU83U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U83U12(tU83U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U83U13(tU83U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U83U14(tU83U14Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U83U15(tU83U15Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U83U16(tU83U16Out,~counter[1],~counter[3],counter[4],counter[5]);
and U83U17(tU83U17Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U83U18(tU83U18Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U83U19(tU83U19Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U83U110(tU83U110Out,~counter[4],~counter[5],counter[6]);
and U83U111(tU83U111Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U83U112(tU83U112Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U83U113(tU83U113Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U83U114(tU83U114Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U83U115(tU83U115Out,~counter[0],~counter[2],~counter[3],~counter[5],counter[6]);
and U83U116(tU83U116Out,~counter[0],counter[2],counter[3],counter[5]);
and U83U117(tU83U117Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U83U118(tU83U118Out,counter[0],~counter[2],~counter[3],counter[4],counter[6]);
and U83U119(tU83U119Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U83U120(tU83U120Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:84====================
wire tU84U122Out;
wire tU84U121Out;
wire tU84U131Out;
wire tU84U112Out;
wire tU84U10Out;
wire tU84U117Out;
wire tU84U12Out;
wire tU84U118Out;
wire tU84U110Out;
wire tU84U11Out;
wire tU84U111Out;
wire tU84U126Out;
wire tU84U17Out;
wire tU84U19Out;
wire tU84U116Out;
wire tU84U130Out;
wire tU84U18Out;
wire tU84U123Out;
wire tU84U124Out;
wire tU84U127Out;
wire tU84U119Out;
wire tU84U129Out;
wire tU84U113Out;
wire tU84U13Out;
wire tU84U125Out;
wire tU84U128Out;
wire tU84U15Out;
wire tU84U115Out;
wire tU84U136Out;
wire tU84U114Out;
wire tU84U00Out;
wire tU84U132Out;
wire tU84U135Out;
wire tU84U133Out;
wire tU84U16Out;
wire tU84U120Out;
wire tU84U137Out;
wire tU84U134Out;
wire tU84U14Out;
or U84U00(tU84U00Out,tU84U10Out,tU84U11Out,tU84U12Out,tU84U13Out,tU84U14Out,tU84U15Out,tU84U16Out,tU84U17Out,tU84U18Out,tU84U19Out,tU84U110Out,tU84U111Out,tU84U112Out,tU84U113Out,tU84U114Out,tU84U115Out,tU84U116Out,tU84U117Out,tU84U118Out,tU84U119Out,tU84U120Out,tU84U121Out,tU84U122Out,tU84U123Out,tU84U124Out,tU84U125Out,tU84U126Out,tU84U127Out,tU84U128Out,tU84U129Out,tU84U130Out,tU84U131Out,tU84U132Out,tU84U133Out,tU84U134Out,tU84U135Out,tU84U136Out,tU84U137Out);
and U84U10(tU84U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U84U11(tU84U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U84U12(tU84U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U84U13(tU84U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U84U14(tU84U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U84U15(tU84U15Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U84U16(tU84U16Out,counter[1],~counter[2],counter[4],counter[5]);
and U84U17(tU84U17Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U84U18(tU84U18Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U84U19(tU84U19Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U84U110(tU84U110Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U84U111(tU84U111Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U84U112(tU84U112Out,~counter[1],~counter[3],counter[4],counter[5]);
and U84U113(tU84U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U84U114(tU84U114Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U84U115(tU84U115Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U84U116(tU84U116Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U84U117(tU84U117Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U84U118(tU84U118Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U84U119(tU84U119Out,~counter[4],~counter[5],counter[6]);
and U84U120(tU84U120Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U84U121(tU84U121Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U84U122(tU84U122Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U84U123(tU84U123Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U84U124(tU84U124Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U84U125(tU84U125Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U84U126(tU84U126Out,~counter[0],~counter[2],~counter[3],~counter[5],counter[6]);
and U84U127(tU84U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[5]);
and U84U128(tU84U128Out,~counter[0],counter[2],counter[3],counter[5]);
and U84U129(tU84U129Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U84U130(tU84U130Out,counter[0],~counter[2],~counter[3],counter[4],counter[6]);
and U84U131(tU84U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U84U132(tU84U132Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U84U133(tU84U133Out,~counter[1],counter[2],counter[3],counter[5]);
and U84U134(tU84U134Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U84U135(tU84U135Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U84U136(tU84U136Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U84U137(tU84U137Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:85====================
wire tU85U13Out;
wire tU85U17Out;
wire tU85U18Out;
wire tU85U19Out;
wire tU85U110Out;
wire tU85U00Out;
wire tU85U15Out;
wire tU85U14Out;
wire tU85U16Out;
wire tU85U12Out;
wire tU85U111Out;
wire tU85U112Out;
wire tU85U11Out;
wire tU85U10Out;
or U85U00(tU85U00Out,tU85U10Out,tU85U11Out,tU85U12Out,tU85U13Out,tU85U14Out,tU85U15Out,tU85U16Out,tU85U17Out,tU85U18Out,tU85U19Out,tU85U110Out,tU85U111Out,tU85U112Out);
and U85U10(tU85U10Out,~counter[1],~counter[3],counter[4],counter[6]);
and U85U11(tU85U11Out,counter[1],~counter[2],counter[4],counter[5]);
and U85U12(tU85U12Out,~counter[1],~counter[3],counter[4],counter[5]);
and U85U13(tU85U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U85U14(tU85U14Out,~counter[4],~counter[5],counter[6]);
and U85U15(tU85U15Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U85U16(tU85U16Out,~counter[0],~counter[2],~counter[3],~counter[5],counter[6]);
and U85U17(tU85U17Out,~counter[0],counter[2],counter[3],counter[5]);
and U85U18(tU85U18Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U85U19(tU85U19Out,counter[0],~counter[2],~counter[3],counter[4],counter[6]);
and U85U110(tU85U110Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U85U111(tU85U111Out,~counter[1],counter[2],counter[3],counter[5]);
and U85U112(tU85U112Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:86====================
wire tU86U19Out;
wire tU86U10Out;
wire tU86U125Out;
wire tU86U17Out;
wire tU86U113Out;
wire tU86U124Out;
wire tU86U16Out;
wire tU86U115Out;
wire tU86U123Out;
wire tU86U00Out;
wire tU86U119Out;
wire tU86U11Out;
wire tU86U14Out;
wire tU86U18Out;
wire tU86U120Out;
wire tU86U12Out;
wire tU86U110Out;
wire tU86U116Out;
wire tU86U117Out;
wire tU86U111Out;
wire tU86U15Out;
wire tU86U126Out;
wire tU86U118Out;
wire tU86U122Out;
wire tU86U121Out;
wire tU86U114Out;
wire tU86U13Out;
wire tU86U112Out;
or U86U00(tU86U00Out,tU86U10Out,tU86U11Out,tU86U12Out,tU86U13Out,tU86U14Out,tU86U15Out,tU86U16Out,tU86U17Out,tU86U18Out,tU86U19Out,tU86U110Out,tU86U111Out,tU86U112Out,tU86U113Out,tU86U114Out,tU86U115Out,tU86U116Out,tU86U117Out,tU86U118Out,tU86U119Out,tU86U120Out,tU86U121Out,tU86U122Out,tU86U123Out,tU86U124Out,tU86U125Out,tU86U126Out);
and U86U10(tU86U10Out,~counter[1],~counter[3],counter[4],counter[6]);
and U86U11(tU86U11Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U86U12(tU86U12Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U86U13(tU86U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U86U14(tU86U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U86U15(tU86U15Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U86U16(tU86U16Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U86U17(tU86U17Out,~counter[1],~counter[3],counter[4],counter[5]);
and U86U18(tU86U18Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U86U19(tU86U19Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U86U110(tU86U110Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U86U111(tU86U111Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U86U112(tU86U112Out,~counter[4],~counter[5],counter[6]);
and U86U113(tU86U113Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U86U114(tU86U114Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U86U115(tU86U115Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U86U116(tU86U116Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U86U117(tU86U117Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U86U118(tU86U118Out,~counter[0],counter[2],counter[3],counter[5]);
and U86U119(tU86U119Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U86U120(tU86U120Out,counter[0],~counter[2],~counter[3],counter[4],counter[6]);
and U86U121(tU86U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U86U122(tU86U122Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U86U123(tU86U123Out,~counter[1],counter[2],counter[3],counter[5]);
and U86U124(tU86U124Out,~counter[0],~counter[3],~counter[5],counter[6]);
and U86U125(tU86U125Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U86U126(tU86U126Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:87====================
wire tU87U11Out;
wire tU87U121Out;
wire tU87U111Out;
wire tU87U118Out;
wire tU87U12Out;
wire tU87U119Out;
wire tU87U13Out;
wire tU87U10Out;
wire tU87U15Out;
wire tU87U16Out;
wire tU87U18Out;
wire tU87U19Out;
wire tU87U112Out;
wire tU87U17Out;
wire tU87U114Out;
wire tU87U117Out;
wire tU87U115Out;
wire tU87U00Out;
wire tU87U116Out;
wire tU87U113Out;
wire tU87U110Out;
wire tU87U120Out;
wire tU87U14Out;
or U87U00(tU87U00Out,tU87U10Out,tU87U11Out,tU87U12Out,tU87U13Out,tU87U14Out,tU87U15Out,tU87U16Out,tU87U17Out,tU87U18Out,tU87U19Out,tU87U110Out,tU87U111Out,tU87U112Out,tU87U113Out,tU87U114Out,tU87U115Out,tU87U116Out,tU87U117Out,tU87U118Out,tU87U119Out,tU87U120Out,tU87U121Out);
and U87U10(tU87U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U87U11(tU87U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U87U12(tU87U12Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U87U13(tU87U13Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U87U14(tU87U14Out,counter[1],~counter[2],counter[4],counter[5]);
and U87U15(tU87U15Out,~counter[3],~counter[5],counter[6]);
and U87U16(tU87U16Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U87U17(tU87U17Out,~counter[1],~counter[3],counter[4],counter[5]);
and U87U18(tU87U18Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U87U19(tU87U19Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U87U110(tU87U110Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U87U111(tU87U111Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U87U112(tU87U112Out,~counter[4],~counter[5],counter[6]);
and U87U113(tU87U113Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U87U114(tU87U114Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U87U115(tU87U115Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U87U116(tU87U116Out,~counter[0],counter[2],counter[3],counter[5]);
and U87U117(tU87U117Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U87U118(tU87U118Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U87U119(tU87U119Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U87U120(tU87U120Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U87U121(tU87U121Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:88====================
wire tU88U111Out;
wire tU88U137Out;
wire tU88U142Out;
wire tU88U117Out;
wire tU88U131Out;
wire tU88U125Out;
wire tU88U12Out;
wire tU88U128Out;
wire tU88U14Out;
wire tU88U18Out;
wire tU88U122Out;
wire tU88U132Out;
wire tU88U135Out;
wire tU88U136Out;
wire tU88U120Out;
wire tU88U146Out;
wire tU88U126Out;
wire tU88U134Out;
wire tU88U140Out;
wire tU88U121Out;
wire tU88U15Out;
wire tU88U145Out;
wire tU88U00Out;
wire tU88U16Out;
wire tU88U113Out;
wire tU88U130Out;
wire tU88U133Out;
wire tU88U118Out;
wire tU88U10Out;
wire tU88U129Out;
wire tU88U116Out;
wire tU88U144Out;
wire tU88U138Out;
wire tU88U143Out;
wire tU88U112Out;
wire tU88U139Out;
wire tU88U13Out;
wire tU88U114Out;
wire tU88U110Out;
wire tU88U17Out;
wire tU88U124Out;
wire tU88U127Out;
wire tU88U141Out;
wire tU88U123Out;
wire tU88U19Out;
wire tU88U147Out;
wire tU88U115Out;
wire tU88U119Out;
wire tU88U11Out;
or U88U00(tU88U00Out,tU88U10Out,tU88U11Out,tU88U12Out,tU88U13Out,tU88U14Out,tU88U15Out,tU88U16Out,tU88U17Out,tU88U18Out,tU88U19Out,tU88U110Out,tU88U111Out,tU88U112Out,tU88U113Out,tU88U114Out,tU88U115Out,tU88U116Out,tU88U117Out,tU88U118Out,tU88U119Out,tU88U120Out,tU88U121Out,tU88U122Out,tU88U123Out,tU88U124Out,tU88U125Out,tU88U126Out,tU88U127Out,tU88U128Out,tU88U129Out,tU88U130Out,tU88U131Out,tU88U132Out,tU88U133Out,tU88U134Out,tU88U135Out,tU88U136Out,tU88U137Out,tU88U138Out,tU88U139Out,tU88U140Out,tU88U141Out,tU88U142Out,tU88U143Out,tU88U144Out,tU88U145Out,tU88U146Out,tU88U147Out);
and U88U10(tU88U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U88U11(tU88U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U88U12(tU88U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U88U13(tU88U13Out,~counter[0],~counter[1],~counter[2],~counter[5],counter[6]);
and U88U14(tU88U14Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U88U15(tU88U15Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U88U16(tU88U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U88U17(tU88U17Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U88U18(tU88U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U88U19(tU88U19Out,counter[1],~counter[2],counter[4],counter[5]);
and U88U110(tU88U110Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U88U111(tU88U111Out,~counter[3],~counter[5],counter[6]);
and U88U112(tU88U112Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U88U113(tU88U113Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U88U114(tU88U114Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U88U115(tU88U115Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U88U116(tU88U116Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U88U117(tU88U117Out,~counter[1],~counter[3],counter[4],counter[5]);
and U88U118(tU88U118Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U88U119(tU88U119Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U88U120(tU88U120Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U88U121(tU88U121Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U88U122(tU88U122Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U88U123(tU88U123Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U88U124(tU88U124Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U88U125(tU88U125Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U88U126(tU88U126Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U88U127(tU88U127Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U88U128(tU88U128Out,~counter[4],~counter[5],counter[6]);
and U88U129(tU88U129Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U88U130(tU88U130Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U88U131(tU88U131Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U88U132(tU88U132Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U88U133(tU88U133Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U88U134(tU88U134Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U88U135(tU88U135Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U88U136(tU88U136Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U88U137(tU88U137Out,~counter[0],counter[2],counter[3],counter[5]);
and U88U138(tU88U138Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U88U139(tU88U139Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U88U140(tU88U140Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U88U141(tU88U141Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U88U142(tU88U142Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U88U143(tU88U143Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U88U144(tU88U144Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U88U145(tU88U145Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U88U146(tU88U146Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U88U147(tU88U147Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:89====================
wire tU89U10Out;
wire tU89U00Out;
wire tU89U115Out;
wire tU89U14Out;
wire tU89U113Out;
wire tU89U112Out;
wire tU89U117Out;
wire tU89U123Out;
wire tU89U12Out;
wire tU89U121Out;
wire tU89U111Out;
wire tU89U13Out;
wire tU89U15Out;
wire tU89U125Out;
wire tU89U120Out;
wire tU89U124Out;
wire tU89U19Out;
wire tU89U110Out;
wire tU89U16Out;
wire tU89U18Out;
wire tU89U17Out;
wire tU89U118Out;
wire tU89U116Out;
wire tU89U119Out;
wire tU89U122Out;
wire tU89U127Out;
wire tU89U126Out;
wire tU89U11Out;
wire tU89U114Out;
or U89U00(tU89U00Out,tU89U10Out,tU89U11Out,tU89U12Out,tU89U13Out,tU89U14Out,tU89U15Out,tU89U16Out,tU89U17Out,tU89U18Out,tU89U19Out,tU89U110Out,tU89U111Out,tU89U112Out,tU89U113Out,tU89U114Out,tU89U115Out,tU89U116Out,tU89U117Out,tU89U118Out,tU89U119Out,tU89U120Out,tU89U121Out,tU89U122Out,tU89U123Out,tU89U124Out,tU89U125Out,tU89U126Out,tU89U127Out);
and U89U10(tU89U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U89U11(tU89U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U89U12(tU89U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U89U13(tU89U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U89U14(tU89U14Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U89U15(tU89U15Out,counter[1],~counter[2],counter[4],counter[5]);
and U89U16(tU89U16Out,~counter[3],~counter[5],counter[6]);
and U89U17(tU89U17Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U89U18(tU89U18Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U89U19(tU89U19Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U89U110(tU89U110Out,~counter[1],~counter[3],counter[4],counter[5]);
and U89U111(tU89U111Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U89U112(tU89U112Out,~counter[1],~counter[2],counter[3],counter[4],counter[6]);
and U89U113(tU89U113Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U89U114(tU89U114Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U89U115(tU89U115Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U89U116(tU89U116Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U89U117(tU89U117Out,~counter[4],~counter[5],counter[6]);
and U89U118(tU89U118Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U89U119(tU89U119Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U89U120(tU89U120Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U89U121(tU89U121Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U89U122(tU89U122Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U89U123(tU89U123Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U89U124(tU89U124Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U89U125(tU89U125Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U89U126(tU89U126Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U89U127(tU89U127Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:90====================
wire tU90U128Out;
wire tU90U118Out;
wire tU90U111Out;
wire tU90U125Out;
wire tU90U132Out;
wire tU90U13Out;
wire tU90U134Out;
wire tU90U126Out;
wire tU90U143Out;
wire tU90U124Out;
wire tU90U117Out;
wire tU90U130Out;
wire tU90U114Out;
wire tU90U137Out;
wire tU90U141Out;
wire tU90U136Out;
wire tU90U00Out;
wire tU90U119Out;
wire tU90U17Out;
wire tU90U123Out;
wire tU90U11Out;
wire tU90U120Out;
wire tU90U127Out;
wire tU90U10Out;
wire tU90U139Out;
wire tU90U112Out;
wire tU90U18Out;
wire tU90U133Out;
wire tU90U15Out;
wire tU90U14Out;
wire tU90U12Out;
wire tU90U121Out;
wire tU90U138Out;
wire tU90U135Out;
wire tU90U122Out;
wire tU90U115Out;
wire tU90U129Out;
wire tU90U110Out;
wire tU90U16Out;
wire tU90U142Out;
wire tU90U140Out;
wire tU90U144Out;
wire tU90U113Out;
wire tU90U131Out;
wire tU90U19Out;
wire tU90U116Out;
or U90U00(tU90U00Out,tU90U10Out,tU90U11Out,tU90U12Out,tU90U13Out,tU90U14Out,tU90U15Out,tU90U16Out,tU90U17Out,tU90U18Out,tU90U19Out,tU90U110Out,tU90U111Out,tU90U112Out,tU90U113Out,tU90U114Out,tU90U115Out,tU90U116Out,tU90U117Out,tU90U118Out,tU90U119Out,tU90U120Out,tU90U121Out,tU90U122Out,tU90U123Out,tU90U124Out,tU90U125Out,tU90U126Out,tU90U127Out,tU90U128Out,tU90U129Out,tU90U130Out,tU90U131Out,tU90U132Out,tU90U133Out,tU90U134Out,tU90U135Out,tU90U136Out,tU90U137Out,tU90U138Out,tU90U139Out,tU90U140Out,tU90U141Out,tU90U142Out,tU90U143Out,tU90U144Out);
and U90U10(tU90U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U90U11(tU90U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U90U12(tU90U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U90U13(tU90U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U90U14(tU90U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U90U15(tU90U15Out,~counter[0],~counter[2],~counter[5],counter[6]);
and U90U16(tU90U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U90U17(tU90U17Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U90U18(tU90U18Out,counter[1],~counter[2],counter[4],counter[5]);
and U90U19(tU90U19Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U90U110(tU90U110Out,~counter[3],~counter[5],counter[6]);
and U90U111(tU90U111Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U90U112(tU90U112Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U90U113(tU90U113Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U90U114(tU90U114Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U90U115(tU90U115Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U90U116(tU90U116Out,~counter[1],~counter[3],counter[4],counter[5]);
and U90U117(tU90U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U90U118(tU90U118Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U90U119(tU90U119Out,~counter[1],~counter[2],counter[3],counter[4],counter[6]);
and U90U120(tU90U120Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U90U121(tU90U121Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U90U122(tU90U122Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U90U123(tU90U123Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U90U124(tU90U124Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U90U125(tU90U125Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U90U126(tU90U126Out,~counter[4],~counter[5],counter[6]);
and U90U127(tU90U127Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U90U128(tU90U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U90U129(tU90U129Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U90U130(tU90U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U90U131(tU90U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U90U132(tU90U132Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U90U133(tU90U133Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U90U134(tU90U134Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U90U135(tU90U135Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U90U136(tU90U136Out,~counter[0],counter[2],counter[3],counter[5]);
and U90U137(tU90U137Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U90U138(tU90U138Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U90U139(tU90U139Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U90U140(tU90U140Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U90U141(tU90U141Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U90U142(tU90U142Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U90U143(tU90U143Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U90U144(tU90U144Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:91====================
wire tU91U110Out;
wire tU91U126Out;
wire tU91U19Out;
wire tU91U11Out;
wire tU91U118Out;
wire tU91U17Out;
wire tU91U113Out;
wire tU91U111Out;
wire tU91U13Out;
wire tU91U121Out;
wire tU91U119Out;
wire tU91U122Out;
wire tU91U00Out;
wire tU91U12Out;
wire tU91U116Out;
wire tU91U120Out;
wire tU91U124Out;
wire tU91U15Out;
wire tU91U112Out;
wire tU91U18Out;
wire tU91U14Out;
wire tU91U115Out;
wire tU91U125Out;
wire tU91U117Out;
wire tU91U123Out;
wire tU91U10Out;
wire tU91U114Out;
wire tU91U16Out;
or U91U00(tU91U00Out,tU91U10Out,tU91U11Out,tU91U12Out,tU91U13Out,tU91U14Out,tU91U15Out,tU91U16Out,tU91U17Out,tU91U18Out,tU91U19Out,tU91U110Out,tU91U111Out,tU91U112Out,tU91U113Out,tU91U114Out,tU91U115Out,tU91U116Out,tU91U117Out,tU91U118Out,tU91U119Out,tU91U120Out,tU91U121Out,tU91U122Out,tU91U123Out,tU91U124Out,tU91U125Out,tU91U126Out);
and U91U10(tU91U10Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U91U11(tU91U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U91U12(tU91U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U91U13(tU91U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U91U14(tU91U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U91U15(tU91U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U91U16(tU91U16Out,counter[1],~counter[2],counter[4],counter[5]);
and U91U17(tU91U17Out,~counter[3],~counter[5],counter[6]);
and U91U18(tU91U18Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U91U19(tU91U19Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U91U110(tU91U110Out,~counter[1],~counter[3],counter[4],counter[5]);
and U91U111(tU91U111Out,~counter[1],~counter[2],counter[3],counter[4],counter[6]);
and U91U112(tU91U112Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U91U113(tU91U113Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U91U114(tU91U114Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U91U115(tU91U115Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U91U116(tU91U116Out,~counter[4],~counter[5],counter[6]);
and U91U117(tU91U117Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U91U118(tU91U118Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U91U119(tU91U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U91U120(tU91U120Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U91U121(tU91U121Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U91U122(tU91U122Out,counter[1],~counter[2],counter[4],counter[6]);
and U91U123(tU91U123Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U91U124(tU91U124Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U91U125(tU91U125Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U91U126(tU91U126Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:92====================
wire tU92U13Out;
wire tU92U110Out;
wire tU92U17Out;
wire tU92U00Out;
wire tU92U19Out;
wire tU92U120Out;
wire tU92U119Out;
wire tU92U116Out;
wire tU92U14Out;
wire tU92U123Out;
wire tU92U11Out;
wire tU92U115Out;
wire tU92U122Out;
wire tU92U112Out;
wire tU92U15Out;
wire tU92U10Out;
wire tU92U125Out;
wire tU92U111Out;
wire tU92U114Out;
wire tU92U113Out;
wire tU92U16Out;
wire tU92U12Out;
wire tU92U118Out;
wire tU92U124Out;
wire tU92U18Out;
wire tU92U121Out;
wire tU92U117Out;
or U92U00(tU92U00Out,tU92U10Out,tU92U11Out,tU92U12Out,tU92U13Out,tU92U14Out,tU92U15Out,tU92U16Out,tU92U17Out,tU92U18Out,tU92U19Out,tU92U110Out,tU92U111Out,tU92U112Out,tU92U113Out,tU92U114Out,tU92U115Out,tU92U116Out,tU92U117Out,tU92U118Out,tU92U119Out,tU92U120Out,tU92U121Out,tU92U122Out,tU92U123Out,tU92U124Out,tU92U125Out);
and U92U10(tU92U10Out,~counter[0],~counter[1],counter[4],counter[6]);
and U92U11(tU92U11Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U92U12(tU92U12Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U92U13(tU92U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U92U14(tU92U14Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U92U15(tU92U15Out,~counter[3],~counter[5],counter[6]);
and U92U16(tU92U16Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U92U17(tU92U17Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U92U18(tU92U18Out,~counter[1],~counter[3],counter[4],counter[5]);
and U92U19(tU92U19Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U92U110(tU92U110Out,~counter[1],~counter[2],counter[3],counter[4],counter[6]);
and U92U111(tU92U111Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U92U112(tU92U112Out,~counter[4],~counter[5],counter[6]);
and U92U113(tU92U113Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U92U114(tU92U114Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U92U115(tU92U115Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U92U116(tU92U116Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U92U117(tU92U117Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U92U118(tU92U118Out,~counter[0],counter[2],counter[3],counter[5]);
and U92U119(tU92U119Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U92U120(tU92U120Out,counter[1],~counter[2],counter[4],counter[6]);
and U92U121(tU92U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U92U122(tU92U122Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U92U123(tU92U123Out,~counter[1],counter[2],counter[3],counter[5]);
and U92U124(tU92U124Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U92U125(tU92U125Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:93====================
wire tU93U14Out;
wire tU93U18Out;
wire tU93U00Out;
wire tU93U15Out;
wire tU93U10Out;
wire tU93U19Out;
wire tU93U11Out;
wire tU93U16Out;
wire tU93U13Out;
wire tU93U12Out;
wire tU93U17Out;
or U93U00(tU93U00Out,tU93U10Out,tU93U11Out,tU93U12Out,tU93U13Out,tU93U14Out,tU93U15Out,tU93U16Out,tU93U17Out,tU93U18Out,tU93U19Out);
and U93U10(tU93U10Out,counter[1],~counter[2],counter[4],counter[5]);
and U93U11(tU93U11Out,~counter[3],~counter[5],counter[6]);
and U93U12(tU93U12Out,~counter[1],~counter[3],counter[4],counter[5]);
and U93U13(tU93U13Out,~counter[4],~counter[5],counter[6]);
and U93U14(tU93U14Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U93U15(tU93U15Out,~counter[1],~counter[5],counter[6]);
and U93U16(tU93U16Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U93U17(tU93U17Out,counter[1],~counter[2],counter[4],counter[6]);
and U93U18(tU93U18Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U93U19(tU93U19Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:94====================
wire tU94U13Out;
wire tU94U14Out;
wire tU94U16Out;
wire tU94U18Out;
wire tU94U120Out;
wire tU94U124Out;
wire tU94U17Out;
wire tU94U136Out;
wire tU94U114Out;
wire tU94U123Out;
wire tU94U137Out;
wire tU94U126Out;
wire tU94U110Out;
wire tU94U112Out;
wire tU94U128Out;
wire tU94U118Out;
wire tU94U113Out;
wire tU94U15Out;
wire tU94U117Out;
wire tU94U121Out;
wire tU94U134Out;
wire tU94U111Out;
wire tU94U116Out;
wire tU94U12Out;
wire tU94U11Out;
wire tU94U131Out;
wire tU94U00Out;
wire tU94U127Out;
wire tU94U10Out;
wire tU94U115Out;
wire tU94U135Out;
wire tU94U132Out;
wire tU94U129Out;
wire tU94U122Out;
wire tU94U138Out;
wire tU94U119Out;
wire tU94U130Out;
wire tU94U133Out;
wire tU94U19Out;
wire tU94U125Out;
or U94U00(tU94U00Out,tU94U10Out,tU94U11Out,tU94U12Out,tU94U13Out,tU94U14Out,tU94U15Out,tU94U16Out,tU94U17Out,tU94U18Out,tU94U19Out,tU94U110Out,tU94U111Out,tU94U112Out,tU94U113Out,tU94U114Out,tU94U115Out,tU94U116Out,tU94U117Out,tU94U118Out,tU94U119Out,tU94U120Out,tU94U121Out,tU94U122Out,tU94U123Out,tU94U124Out,tU94U125Out,tU94U126Out,tU94U127Out,tU94U128Out,tU94U129Out,tU94U130Out,tU94U131Out,tU94U132Out,tU94U133Out,tU94U134Out,tU94U135Out,tU94U136Out,tU94U137Out,tU94U138Out);
and U94U10(tU94U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U94U11(tU94U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U94U12(tU94U12Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U94U13(tU94U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U94U14(tU94U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U94U15(tU94U15Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U94U16(tU94U16Out,~counter[0],~counter[5],counter[6]);
and U94U17(tU94U17Out,counter[1],~counter[2],counter[4],counter[5]);
and U94U18(tU94U18Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U94U19(tU94U19Out,~counter[3],~counter[5],counter[6]);
and U94U110(tU94U110Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U94U111(tU94U111Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U94U112(tU94U112Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U94U113(tU94U113Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U94U114(tU94U114Out,~counter[1],~counter[3],counter[4],counter[5]);
and U94U115(tU94U115Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U94U116(tU94U116Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U94U117(tU94U117Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U94U118(tU94U118Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U94U119(tU94U119Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U94U120(tU94U120Out,~counter[4],~counter[5],counter[6]);
and U94U121(tU94U121Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U94U122(tU94U122Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U94U123(tU94U123Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U94U124(tU94U124Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U94U125(tU94U125Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U94U126(tU94U126Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U94U127(tU94U127Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U94U128(tU94U128Out,~counter[1],~counter[5],counter[6]);
and U94U129(tU94U129Out,~counter[0],counter[2],counter[3],counter[5]);
and U94U130(tU94U130Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U94U131(tU94U131Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U94U132(tU94U132Out,counter[1],~counter[2],counter[4],counter[6]);
and U94U133(tU94U133Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U94U134(tU94U134Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U94U135(tU94U135Out,~counter[1],counter[2],counter[3],counter[5]);
and U94U136(tU94U136Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U94U137(tU94U137Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U94U138(tU94U138Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:95====================
wire tU95U117Out;
wire tU95U110Out;
wire tU95U116Out;
wire tU95U12Out;
wire tU95U119Out;
wire tU95U00Out;
wire tU95U11Out;
wire tU95U118Out;
wire tU95U112Out;
wire tU95U114Out;
wire tU95U111Out;
wire tU95U15Out;
wire tU95U113Out;
wire tU95U18Out;
wire tU95U17Out;
wire tU95U115Out;
wire tU95U10Out;
wire tU95U16Out;
wire tU95U14Out;
wire tU95U120Out;
wire tU95U19Out;
wire tU95U13Out;
or U95U00(tU95U00Out,tU95U10Out,tU95U11Out,tU95U12Out,tU95U13Out,tU95U14Out,tU95U15Out,tU95U16Out,tU95U17Out,tU95U18Out,tU95U19Out,tU95U110Out,tU95U111Out,tU95U112Out,tU95U113Out,tU95U114Out,tU95U115Out,tU95U116Out,tU95U117Out,tU95U118Out,tU95U119Out,tU95U120Out);
and U95U10(tU95U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U95U11(tU95U11Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U95U12(tU95U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U95U13(tU95U13Out,counter[2],counter[4],counter[6]);
and U95U14(tU95U14Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U95U15(tU95U15Out,counter[1],~counter[2],counter[4],counter[5]);
and U95U16(tU95U16Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U95U17(tU95U17Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U95U18(tU95U18Out,~counter[1],~counter[3],counter[4],counter[5]);
and U95U19(tU95U19Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U95U110(tU95U110Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U95U111(tU95U111Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U95U112(tU95U112Out,~counter[4],~counter[5],counter[6]);
and U95U113(tU95U113Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U95U114(tU95U114Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U95U115(tU95U115Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U95U116(tU95U116Out,~counter[1],~counter[5],counter[6]);
and U95U117(tU95U117Out,counter[1],~counter[2],counter[4],counter[6]);
and U95U118(tU95U118Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U95U119(tU95U119Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U95U120(tU95U120Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:96====================
wire tU96U120Out;
wire tU96U11Out;
wire tU96U116Out;
wire tU96U16Out;
wire tU96U123Out;
wire tU96U115Out;
wire tU96U147Out;
wire tU96U129Out;
wire tU96U18Out;
wire tU96U128Out;
wire tU96U121Out;
wire tU96U136Out;
wire tU96U14Out;
wire tU96U19Out;
wire tU96U113Out;
wire tU96U119Out;
wire tU96U144Out;
wire tU96U125Out;
wire tU96U111Out;
wire tU96U117Out;
wire tU96U134Out;
wire tU96U142Out;
wire tU96U112Out;
wire tU96U122Out;
wire tU96U135Out;
wire tU96U133Out;
wire tU96U141Out;
wire tU96U12Out;
wire tU96U127Out;
wire tU96U140Out;
wire tU96U00Out;
wire tU96U118Out;
wire tU96U146Out;
wire tU96U10Out;
wire tU96U139Out;
wire tU96U149Out;
wire tU96U148Out;
wire tU96U132Out;
wire tU96U131Out;
wire tU96U13Out;
wire tU96U15Out;
wire tU96U17Out;
wire tU96U145Out;
wire tU96U138Out;
wire tU96U130Out;
wire tU96U110Out;
wire tU96U124Out;
wire tU96U114Out;
wire tU96U137Out;
wire tU96U143Out;
wire tU96U126Out;
or U96U00(tU96U00Out,tU96U10Out,tU96U11Out,tU96U12Out,tU96U13Out,tU96U14Out,tU96U15Out,tU96U16Out,tU96U17Out,tU96U18Out,tU96U19Out,tU96U110Out,tU96U111Out,tU96U112Out,tU96U113Out,tU96U114Out,tU96U115Out,tU96U116Out,tU96U117Out,tU96U118Out,tU96U119Out,tU96U120Out,tU96U121Out,tU96U122Out,tU96U123Out,tU96U124Out,tU96U125Out,tU96U126Out,tU96U127Out,tU96U128Out,tU96U129Out,tU96U130Out,tU96U131Out,tU96U132Out,tU96U133Out,tU96U134Out,tU96U135Out,tU96U136Out,tU96U137Out,tU96U138Out,tU96U139Out,tU96U140Out,tU96U141Out,tU96U142Out,tU96U143Out,tU96U144Out,tU96U145Out,tU96U146Out,tU96U147Out,tU96U148Out,tU96U149Out);
and U96U10(tU96U10Out,counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U96U11(tU96U11Out,counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U96U12(tU96U12Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U96U13(tU96U13Out,~counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[6]);
and U96U14(tU96U14Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U96U15(tU96U15Out,counter[2],counter[4],counter[6]);
and U96U16(tU96U16Out,counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U96U17(tU96U17Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U96U18(tU96U18Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U96U19(tU96U19Out,counter[1],~counter[2],counter[4],counter[5]);
and U96U110(tU96U110Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U96U111(tU96U111Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U96U112(tU96U112Out,counter[0],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U96U113(tU96U113Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U96U114(tU96U114Out,~counter[0],~counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U96U115(tU96U115Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U96U116(tU96U116Out,~counter[1],~counter[3],counter[4],counter[5]);
and U96U117(tU96U117Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U96U118(tU96U118Out,counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U96U119(tU96U119Out,counter[0],~counter[1],counter[2],counter[3],~counter[4]);
and U96U120(tU96U120Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U96U121(tU96U121Out,~counter[0],counter[2],counter[3],~counter[4],~counter[5]);
and U96U122(tU96U122Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U96U123(tU96U123Out,counter[0],~counter[1],~counter[3],~counter[4],~counter[5],~counter[6]);
and U96U124(tU96U124Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U96U125(tU96U125Out,counter[0],counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U96U126(tU96U126Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U96U127(tU96U127Out,~counter[4],~counter[5],counter[6]);
and U96U128(tU96U128Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[6]);
and U96U129(tU96U129Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U96U130(tU96U130Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U96U131(tU96U131Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U96U132(tU96U132Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U96U133(tU96U133Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U96U134(tU96U134Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U96U135(tU96U135Out,~counter[0],~counter[1],~counter[2],counter[6]);
and U96U136(tU96U136Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U96U137(tU96U137Out,~counter[1],~counter[5],counter[6]);
and U96U138(tU96U138Out,~counter[0],counter[2],counter[3],counter[5]);
and U96U139(tU96U139Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U96U140(tU96U140Out,~counter[0],~counter[1],counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U96U141(tU96U141Out,counter[1],~counter[2],counter[4],counter[6]);
and U96U142(tU96U142Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U96U143(tU96U143Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U96U144(tU96U144Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U96U145(tU96U145Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U96U146(tU96U146Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U96U147(tU96U147Out,~counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U96U148(tU96U148Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
and U96U149(tU96U149Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:97====================
wire tU97U113Out;
wire tU97U110Out;
wire tU97U112Out;
wire tU97U15Out;
wire tU97U00Out;
wire tU97U16Out;
wire tU97U111Out;
wire tU97U14Out;
wire tU97U12Out;
wire tU97U18Out;
wire tU97U11Out;
wire tU97U10Out;
wire tU97U19Out;
wire tU97U17Out;
wire tU97U13Out;
or U97U00(tU97U00Out,tU97U10Out,tU97U11Out,tU97U12Out,tU97U13Out,tU97U14Out,tU97U15Out,tU97U16Out,tU97U17Out,tU97U18Out,tU97U19Out,tU97U110Out,tU97U111Out,tU97U112Out,tU97U113Out);
and U97U10(tU97U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U97U11(tU97U11Out,counter[2],counter[4],counter[6]);
and U97U12(tU97U12Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U97U13(tU97U13Out,counter[1],~counter[2],counter[4],counter[5]);
and U97U14(tU97U14Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U97U15(tU97U15Out,counter[0],~counter[2],~counter[3],counter[4],counter[5]);
and U97U16(tU97U16Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U97U17(tU97U17Out,~counter[4],~counter[5],counter[6]);
and U97U18(tU97U18Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U97U19(tU97U19Out,~counter[1],~counter[2],counter[6]);
and U97U110(tU97U110Out,counter[1],~counter[2],counter[4],counter[6]);
and U97U111(tU97U111Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U97U112(tU97U112Out,~counter[0],~counter[2],counter[3],~counter[4],~counter[5]);
and U97U113(tU97U113Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:98====================
wire tU98U18Out;
wire tU98U12Out;
wire tU98U122Out;
wire tU98U116Out;
wire tU98U112Out;
wire tU98U118Out;
wire tU98U110Out;
wire tU98U115Out;
wire tU98U14Out;
wire tU98U13Out;
wire tU98U11Out;
wire tU98U125Out;
wire tU98U17Out;
wire tU98U124Out;
wire tU98U10Out;
wire tU98U114Out;
wire tU98U123Out;
wire tU98U19Out;
wire tU98U121Out;
wire tU98U111Out;
wire tU98U113Out;
wire tU98U00Out;
wire tU98U16Out;
wire tU98U119Out;
wire tU98U117Out;
wire tU98U15Out;
wire tU98U120Out;
or U98U00(tU98U00Out,tU98U10Out,tU98U11Out,tU98U12Out,tU98U13Out,tU98U14Out,tU98U15Out,tU98U16Out,tU98U17Out,tU98U18Out,tU98U19Out,tU98U110Out,tU98U111Out,tU98U112Out,tU98U113Out,tU98U114Out,tU98U115Out,tU98U116Out,tU98U117Out,tU98U118Out,tU98U119Out,tU98U120Out,tU98U121Out,tU98U122Out,tU98U123Out,tU98U124Out,tU98U125Out);
and U98U10(tU98U10Out,~counter[0],~counter[2],counter[6]);
and U98U11(tU98U11Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U98U12(tU98U12Out,counter[2],counter[4],counter[6]);
and U98U13(tU98U13Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U98U14(tU98U14Out,counter[1],~counter[2],counter[4],counter[5]);
and U98U15(tU98U15Out,counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U98U16(tU98U16Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U98U17(tU98U17Out,~counter[1],~counter[3],counter[4],counter[5]);
and U98U18(tU98U18Out,~counter[0],counter[1],~counter[2],~counter[3],counter[5],~counter[6]);
and U98U19(tU98U19Out,counter[0],~counter[1],~counter[2],~counter[4],~counter[5],~counter[6]);
and U98U110(tU98U110Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U98U111(tU98U111Out,~counter[4],~counter[5],counter[6]);
and U98U112(tU98U112Out,counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U98U113(tU98U113Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U98U114(tU98U114Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U98U115(tU98U115Out,~counter[1],~counter[2],counter[3],counter[4],counter[5]);
and U98U116(tU98U116Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U98U117(tU98U117Out,~counter[1],~counter[2],counter[6]);
and U98U118(tU98U118Out,~counter[0],counter[2],counter[3],counter[5]);
and U98U119(tU98U119Out,counter[0],counter[1],counter[2],counter[3],~counter[4],counter[5]);
and U98U120(tU98U120Out,counter[1],~counter[2],counter[4],counter[6]);
and U98U121(tU98U121Out,~counter[0],counter[1],counter[2],~counter[3],~counter[4],counter[5]);
and U98U122(tU98U122Out,~counter[0],counter[1],~counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U98U123(tU98U123Out,~counter[1],counter[2],counter[3],counter[5]);
and U98U124(tU98U124Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U98U125(tU98U125Out,counter[2],counter[4],counter[5]);

//====================Truthtable Variable:99====================
wire tU99U119Out;
wire tU99U122Out;
wire tU99U115Out;
wire tU99U12Out;
wire tU99U10Out;
wire tU99U15Out;
wire tU99U112Out;
wire tU99U17Out;
wire tU99U116Out;
wire tU99U121Out;
wire tU99U110Out;
wire tU99U111Out;
wire tU99U118Out;
wire tU99U14Out;
wire tU99U117Out;
wire tU99U00Out;
wire tU99U19Out;
wire tU99U13Out;
wire tU99U123Out;
wire tU99U11Out;
wire tU99U16Out;
wire tU99U113Out;
wire tU99U114Out;
wire tU99U18Out;
wire tU99U120Out;
or U99U00(tU99U00Out,tU99U10Out,tU99U11Out,tU99U12Out,tU99U13Out,tU99U14Out,tU99U15Out,tU99U16Out,tU99U17Out,tU99U18Out,tU99U19Out,tU99U110Out,tU99U111Out,tU99U112Out,tU99U113Out,tU99U114Out,tU99U115Out,tU99U116Out,tU99U117Out,tU99U118Out,tU99U119Out,tU99U120Out,tU99U121Out,tU99U122Out,tU99U123Out);
and U99U10(tU99U10Out,counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U99U11(tU99U11Out,counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U99U12(tU99U12Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U99U13(tU99U13Out,counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U99U14(tU99U14Out,~counter[0],~counter[1],counter[3],~counter[4],counter[5]);
and U99U15(tU99U15Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U99U16(tU99U16Out,~counter[0],~counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U99U17(tU99U17Out,~counter[0],~counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U99U18(tU99U18Out,counter[0],~counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U99U19(tU99U19Out,counter[0],counter[3],counter[4],~counter[5],~counter[6]);
and U99U110(tU99U110Out,counter[2],~counter[4],counter[5]);
and U99U111(tU99U111Out,~counter[0],~counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U99U112(tU99U112Out,~counter[0],counter[1],counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U99U113(tU99U113Out,~counter[1],~counter[2],~counter[3],counter[4],counter[5]);
and U99U114(tU99U114Out,~counter[0],counter[1],~counter[2],~counter[3],counter[4],~counter[5],~counter[6]);
and U99U115(tU99U115Out,counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U99U116(tU99U116Out,~counter[0],counter[1],counter[2],counter[3],~counter[4],~counter[5],~counter[6]);
and U99U117(tU99U117Out,counter[0],counter[1],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U99U118(tU99U118Out,~counter[0],counter[1],~counter[2],counter[3],~counter[4],counter[5]);
and U99U119(tU99U119Out,~counter[0],~counter[1],counter[2],~counter[3],~counter[4],~counter[5],~counter[6]);
and U99U120(tU99U120Out,~counter[0],counter[1],~counter[2],counter[3],counter[4],~counter[5],~counter[6]);
and U99U121(tU99U121Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[4],~counter[6]);
and U99U122(tU99U122Out,~counter[0],~counter[2],~counter[3],~counter[4],counter[5],~counter[6]);
and U99U123(tU99U123Out,counter[0],~counter[1],~counter[2],~counter[3],~counter[5],~counter[6]);
//print("assign lamb={%s}"% (''.join([("tU%dU00Out,"%i) for i in range(0,100)])[:-1]))
assign lamb={tU0U00Out,tU1U00Out,tU2U00Out,tU3U00Out,tU4U00Out,tU5U00Out,tU6U00Out,tU7U00Out,tU8U00Out,tU9U00Out,tU10U00Out,tU11U00Out,tU12U00Out,tU13U00Out,tU14U00Out,tU15U00Out,tU16U00Out,tU17U00Out,tU18U00Out,tU19U00Out,tU20U00Out,tU21U00Out,tU22U00Out,tU23U00Out,tU24U00Out,tU25U00Out,tU26U00Out,tU27U00Out,tU28U00Out,tU29U00Out,tU30U00Out,tU31U00Out,tU32U00Out,tU33U00Out,tU34U00Out,tU35U00Out,tU36U00Out,tU37U00Out,tU38U00Out,tU39U00Out,tU40U00Out,tU41U00Out,tU42U00Out,tU43U00Out,tU44U00Out,tU45U00Out,tU46U00Out,tU47U00Out,tU48U00Out,tU49U00Out,tU50U00Out,tU51U00Out,tU52U00Out,tU53U00Out,tU54U00Out,tU55U00Out,tU56U00Out,tU57U00Out,tU58U00Out,tU59U00Out,tU60U00Out,tU61U00Out,tU62U00Out,tU63U00Out,tU64U00Out,tU65U00Out,tU66U00Out,tU67U00Out,tU68U00Out,tU69U00Out,tU70U00Out,tU71U00Out,tU72U00Out,tU73U00Out,tU74U00Out,tU75U00Out,tU76U00Out,tU77U00Out,tU78U00Out,tU79U00Out,tU80U00Out,tU81U00Out,tU82U00Out,tU83U00Out,tU84U00Out,tU85U00Out,tU86U00Out,tU87U00Out,tU88U00Out,tU89U00Out,tU90U00Out,tU91U00Out,tU92U00Out,tU93U00Out,tU94U00Out,tU95U00Out,tU96U00Out,tU97U00Out,tU98U00Out,tU99U00Out};
endmodule


`timescale 1us/1us
module testlamb100Control();
    reg trigger;
    reg sysRst;
    wire [99:0] lamb;
    wire [6:0] counter;
    
    lamb100Control U1(
        trigger,
        sysRst,
        counter,
        lamb
    );
    initial begin
        sysRst<=1;
        trigger<=0;
        #5 sysRst<=0;
        #2
        sysRst<=1;
        #2
        sysRst<=0;
        #12000 $stop;
        
    end
    always begin
        #5
        trigger<=~trigger;
    end


endmodule


