 module lamp100Prom(
    input [9:0]address,
    output reg [15:0]data
);
always@(*) begin
    case(address)
		10'h0:data=16'b1111111111111111;//STATE:1	SEG:1	COUNTER:0	
		10'h1:data=16'b1111111111111111;//STATE:1	SEG:2	COUNTER:1	
		10'h2:data=16'b1111111111111111;//STATE:1	SEG:3	COUNTER:2	
		10'h3:data=16'b1111111111111111;//STATE:1	SEG:4	COUNTER:3	
		10'h4:data=16'b1111111111111111;//STATE:1	SEG:5	COUNTER:4	
		10'h5:data=16'b1111111111111111;//STATE:1	SEG:6	COUNTER:5	
		10'h6:data=16'b1111000000000000;//STATE:1	SEG:7	COUNTER:6	
		10'h7:data=16'b1010101010101010;//STATE:2	SEG:1	COUNTER:7	
		10'h8:data=16'b1010101010101010;//STATE:2	SEG:2	COUNTER:8	
		10'h9:data=16'b1010101010101010;//STATE:2	SEG:3	COUNTER:9	
		10'ha:data=16'b1010101010101010;//STATE:2	SEG:4	COUNTER:10	
		10'hb:data=16'b1010101010101010;//STATE:2	SEG:5	COUNTER:11	
		10'hc:data=16'b1010101010101010;//STATE:2	SEG:6	COUNTER:12	
		10'hd:data=16'b1010000000000000;//STATE:2	SEG:7	COUNTER:13	
		10'he:data=16'b1000111000111000;//STATE:3	SEG:1	COUNTER:14	
		10'hf:data=16'b1110001110001110;//STATE:3	SEG:2	COUNTER:15	
		10'h10:data=16'b0011100011100011;//STATE:3	SEG:3	COUNTER:16	
		10'h11:data=16'b1000111000111000;//STATE:3	SEG:4	COUNTER:17	
		10'h12:data=16'b1110001110001110;//STATE:3	SEG:5	COUNTER:18	
		10'h13:data=16'b0011100011100011;//STATE:3	SEG:6	COUNTER:19	
		10'h14:data=16'b1000000000000000;//STATE:3	SEG:7	COUNTER:20	
		10'h15:data=16'b1001111100101001;//STATE:4	SEG:1	COUNTER:21	
		10'h16:data=16'b1111001010011111;//STATE:4	SEG:2	COUNTER:22	
		10'h17:data=16'b0010100111110010;//STATE:4	SEG:3	COUNTER:23	
		10'h18:data=16'b1001111100101001;//STATE:4	SEG:4	COUNTER:24	
		10'h19:data=16'b1111001010011111;//STATE:4	SEG:5	COUNTER:25	
		10'h1a:data=16'b0010100111110010;//STATE:4	SEG:6	COUNTER:26	
		10'h1b:data=16'b1001000000000000;//STATE:4	SEG:7	COUNTER:27	
		10'h1c:data=16'b1001011101101011;//STATE:5	SEG:1	COUNTER:28	
		10'h1d:data=16'b1110001000011011;//STATE:5	SEG:2	COUNTER:29	
		10'h1e:data=16'b0000100011111010;//STATE:5	SEG:3	COUNTER:30	
		10'h1f:data=16'b1101110100111001;//STATE:5	SEG:4	COUNTER:31	
		10'h20:data=16'b0111011010111110;//STATE:5	SEG:5	COUNTER:32	
		10'h21:data=16'b0010000110110000;//STATE:5	SEG:6	COUNTER:33	
		10'h22:data=16'b1000000000000000;//STATE:5	SEG:7	COUNTER:34	
		10'h23:data=16'b1001001101111011;//STATE:6	SEG:1	COUNTER:35	
		10'h24:data=16'b1010001100011111;//STATE:6	SEG:2	COUNTER:36	
		10'h25:data=16'b0001100010111011;//STATE:6	SEG:3	COUNTER:37	
		10'h26:data=16'b1101100100101001;//STATE:6	SEG:4	COUNTER:38	
		10'h27:data=16'b0011011110111010;//STATE:6	SEG:5	COUNTER:39	
		10'h28:data=16'b0011000111110001;//STATE:6	SEG:6	COUNTER:40	
		10'h29:data=16'b1000000000000000;//STATE:6	SEG:7	COUNTER:41	
		10'h2a:data=16'b1001000101111111;//STATE:7	SEG:1	COUNTER:42	
		10'h2b:data=16'b1010101100001111;//STATE:7	SEG:2	COUNTER:43	
		10'h2c:data=16'b0011100011111011;//STATE:7	SEG:3	COUNTER:44	
		10'h2d:data=16'b0101100000101011;//STATE:7	SEG:4	COUNTER:45	
		10'h2e:data=16'b0011001110110010;//STATE:7	SEG:5	COUNTER:46	
		10'h2f:data=16'b0010000111010001;//STATE:7	SEG:6	COUNTER:47	
		10'h30:data=16'b1100000000000000;//STATE:7	SEG:7	COUNTER:48	
		10'h31:data=16'b1001000001111110;//STATE:8	SEG:1	COUNTER:49	
		10'h32:data=16'b1010101000001110;//STATE:8	SEG:2	COUNTER:50	
		10'h33:data=16'b0011100111111010;//STATE:8	SEG:3	COUNTER:51	
		10'h34:data=16'b0101100100101010;//STATE:8	SEG:4	COUNTER:52	
		10'h35:data=16'b0011001010110011;//STATE:8	SEG:5	COUNTER:53	
		10'h36:data=16'b0010000011010000;//STATE:8	SEG:6	COUNTER:54	
		10'h37:data=16'b1100000000000000;//STATE:8	SEG:7	COUNTER:55	
		10'h38:data=16'b1001000011111110;//STATE:9	SEG:1	COUNTER:56	
		10'h39:data=16'b1110101000101110;//STATE:9	SEG:2	COUNTER:57	
		10'h3a:data=16'b0010100111110010;//STATE:9	SEG:3	COUNTER:58	
		10'h3b:data=16'b0101110100101000;//STATE:9	SEG:4	COUNTER:59	
		10'h3c:data=16'b0011001110110011;//STATE:9	SEG:5	COUNTER:60	
		10'h3d:data=16'b1010000010010000;//STATE:9	SEG:6	COUNTER:61	
		10'h3e:data=16'b1110000000000000;//STATE:9	SEG:7	COUNTER:62	
		10'h3f:data=16'b1001000010111110;//STATE:10	SEG:1	COUNTER:63	
		10'h40:data=16'b1111101000101010;//STATE:10	SEG:2	COUNTER:64	
		10'h41:data=16'b0010100011110010;//STATE:10	SEG:3	COUNTER:65	
		10'h42:data=16'b0001110100111000;//STATE:10	SEG:4	COUNTER:66	
		10'h43:data=16'b0011011110110010;//STATE:10	SEG:5	COUNTER:67	
		10'h44:data=16'b1010000011010000;//STATE:10	SEG:6	COUNTER:68	
		10'h45:data=16'b1111000000000000;//STATE:10	SEG:7	COUNTER:69	
		10'h46:data=16'b1001000010011110;//STATE:11	SEG:1	COUNTER:70	
		10'h47:data=16'b1111111000101010;//STATE:11	SEG:2	COUNTER:71	
		10'h48:data=16'b1010100011100010;//STATE:11	SEG:3	COUNTER:72	
		10'h49:data=16'b0001111100111000;//STATE:11	SEG:4	COUNTER:73	
		10'h4a:data=16'b0111011110111010;//STATE:11	SEG:5	COUNTER:74	
		10'h4b:data=16'b1010000111010000;//STATE:11	SEG:6	COUNTER:75	
		10'h4c:data=16'b1101000000000000;//STATE:11	SEG:7	COUNTER:76	
		10'h4d:data=16'b1001000010001110;//STATE:12	SEG:1	COUNTER:77	
		10'h4e:data=16'b1111111100101010;//STATE:12	SEG:2	COUNTER:78	
		10'h4f:data=16'b1011100011100011;//STATE:12	SEG:3	COUNTER:79	
		10'h50:data=16'b0001111100101000;//STATE:12	SEG:4	COUNTER:80	
		10'h51:data=16'b0111011010111010;//STATE:12	SEG:5	COUNTER:81	
		10'h52:data=16'b1011000111010001;//STATE:12	SEG:6	COUNTER:82	
		10'h53:data=16'b1101000000000000;//STATE:12	SEG:7	COUNTER:83	
		10'h54:data=16'b1001000010000110;//STATE:13	SEG:1	COUNTER:84	
		10'h55:data=16'b1111111101101010;//STATE:13	SEG:2	COUNTER:85	
		10'h56:data=16'b1011101011100011;//STATE:13	SEG:3	COUNTER:86	
		10'h57:data=16'b0000111100101000;//STATE:13	SEG:4	COUNTER:87	
		10'h58:data=16'b1111011010111110;//STATE:13	SEG:5	COUNTER:88	
		10'h59:data=16'b1011000111110001;//STATE:13	SEG:6	COUNTER:89	
		10'h5a:data=16'b1101000000000000;//STATE:13	SEG:7	COUNTER:90	
		10'h5b:data=16'b1001000010000010;//STATE:14	SEG:1	COUNTER:91	
		10'h5c:data=16'b1111111101111010;//STATE:14	SEG:2	COUNTER:92	
		10'h5d:data=16'b1011101010100011;//STATE:14	SEG:3	COUNTER:93	
		10'h5e:data=16'b0000111000101000;//STATE:14	SEG:4	COUNTER:94	
		10'h5f:data=16'b1111001010111110;//STATE:14	SEG:5	COUNTER:95	
		10'h60:data=16'b1010000111110001;//STATE:14	SEG:6	COUNTER:96	
		10'h61:data=16'b1001000000000000;//STATE:14	SEG:7	COUNTER:97	
		10'h62:data=16'b1001000010000000;//STATE:15	SEG:1	COUNTER:98	
		10'h63:data=16'b1111111101111110;//STATE:15	SEG:2	COUNTER:99	
		10'h64:data=16'b1011101010101011;//STATE:15	SEG:3	COUNTER:100	
		10'h65:data=16'b0000111000111000;//STATE:15	SEG:4	COUNTER:101	
		10'h66:data=16'b1111001010011110;//STATE:15	SEG:5	COUNTER:102	
		10'h67:data=16'b1010000110110001;//STATE:15	SEG:6	COUNTER:103	
		10'h68:data=16'b1001000000000000;//STATE:15	SEG:7	COUNTER:104	
		10'h69:data=16'b1001000010000001;//STATE:16	SEG:1	COUNTER:105	
		10'h6a:data=16'b1111111101111111;//STATE:16	SEG:2	COUNTER:106	
		10'h6b:data=16'b1011101010101010;//STATE:16	SEG:3	COUNTER:107	
		10'h6c:data=16'b0000111000111001;//STATE:16	SEG:4	COUNTER:108	
		10'h6d:data=16'b1111001010011111;//STATE:16	SEG:5	COUNTER:109	
		10'h6e:data=16'b1010000110110000;//STATE:16	SEG:6	COUNTER:110	
		10'h6f:data=16'b1001000000000000;//STATE:16	SEG:7	COUNTER:111	
		10'h70:data=16'b1001000010000001;//STATE:17	SEG:1	COUNTER:112	
		10'h71:data=16'b0111111101111111;//STATE:17	SEG:2	COUNTER:113	
		10'h72:data=16'b1111101010101010;//STATE:17	SEG:3	COUNTER:114	
		10'h73:data=16'b0010111000111001;//STATE:17	SEG:4	COUNTER:115	
		10'h74:data=16'b1110001010011111;//STATE:17	SEG:5	COUNTER:116	
		10'h75:data=16'b1010100110110000;//STATE:17	SEG:6	COUNTER:117	
		10'h76:data=16'b1001000000000000;//STATE:17	SEG:7	COUNTER:118	
		10'h77:data=16'b1001000010000001;//STATE:18	SEG:1	COUNTER:119	
		10'h78:data=16'b0011111101111111;//STATE:18	SEG:2	COUNTER:120	
		10'h79:data=16'b1110101010101010;//STATE:18	SEG:3	COUNTER:121	
		10'h7a:data=16'b0010101000111001;//STATE:18	SEG:4	COUNTER:122	
		10'h7b:data=16'b1110001110011111;//STATE:18	SEG:5	COUNTER:123	
		10'h7c:data=16'b1010100111110000;//STATE:18	SEG:6	COUNTER:124	
		10'h7d:data=16'b1001000000000000;//STATE:18	SEG:7	COUNTER:125	
		10'h7e:data=16'b1001000010000001;//STATE:19	SEG:1	COUNTER:126	
		10'h7f:data=16'b0001111101111111;//STATE:19	SEG:2	COUNTER:127	
		10'h80:data=16'b1110111010101010;//STATE:19	SEG:3	COUNTER:128	
		10'h81:data=16'b0010101010111001;//STATE:19	SEG:4	COUNTER:129	
		10'h82:data=16'b1110001110001111;//STATE:19	SEG:5	COUNTER:130	
		10'h83:data=16'b1010100111110010;//STATE:19	SEG:6	COUNTER:131	
		10'h84:data=16'b1001000000000000;//STATE:19	SEG:7	COUNTER:132	
		10'h85:data=16'b1001000010000001;//STATE:20	SEG:1	COUNTER:133	
		10'h86:data=16'b0000111101111111;//STATE:20	SEG:2	COUNTER:134	
		10'h87:data=16'b1110111110101010;//STATE:20	SEG:3	COUNTER:135	
		10'h88:data=16'b0010101010101001;//STATE:20	SEG:4	COUNTER:136	
		10'h89:data=16'b1110001110001110;//STATE:20	SEG:5	COUNTER:137	
		10'h8a:data=16'b1010100111110010;//STATE:20	SEG:6	COUNTER:138	
		10'h8b:data=16'b1000000000000000;//STATE:20	SEG:7	COUNTER:139	
		10'h8c:data=16'b1001000010000001;//STATE:21	SEG:1	COUNTER:140	
		10'h8d:data=16'b0000011101111111;//STATE:21	SEG:2	COUNTER:141	
		10'h8e:data=16'b1110111111101010;//STATE:21	SEG:3	COUNTER:142	
		10'h8f:data=16'b0010101010101011;//STATE:21	SEG:4	COUNTER:143	
		10'h90:data=16'b1110001110001110;//STATE:21	SEG:5	COUNTER:144	
		10'h91:data=16'b1011100111110010;//STATE:21	SEG:6	COUNTER:145	
		10'h92:data=16'b1000000000000000;//STATE:21	SEG:7	COUNTER:146	
		10'h93:data=16'b1001000010000001;//STATE:22	SEG:1	COUNTER:147	
		10'h94:data=16'b0000001101111111;//STATE:22	SEG:2	COUNTER:148	
		10'h95:data=16'b1110111111111010;//STATE:22	SEG:3	COUNTER:149	
		10'h96:data=16'b0010101010101011;//STATE:22	SEG:4	COUNTER:150	
		10'h97:data=16'b1010001110001110;//STATE:22	SEG:5	COUNTER:151	
		10'h98:data=16'b1011100011110010;//STATE:22	SEG:6	COUNTER:152	
		10'h99:data=16'b1000000000000000;//STATE:22	SEG:7	COUNTER:153	
		10'h9a:data=16'b1001000010000001;//STATE:23	SEG:1	COUNTER:154	
		10'h9b:data=16'b0000000101111111;//STATE:23	SEG:2	COUNTER:155	
		10'h9c:data=16'b1110111111111110;//STATE:23	SEG:3	COUNTER:156	
		10'h9d:data=16'b0010101010101011;//STATE:23	SEG:4	COUNTER:157	
		10'h9e:data=16'b1010101110001110;//STATE:23	SEG:5	COUNTER:158	
		10'h9f:data=16'b1011100011100010;//STATE:23	SEG:6	COUNTER:159	
		10'ha0:data=16'b1000000000000000;//STATE:23	SEG:7	COUNTER:160	
		10'ha1:data=16'b1001000010000001;//STATE:24	SEG:1	COUNTER:161	
		10'ha2:data=16'b0000000001111111;//STATE:24	SEG:2	COUNTER:162	
		10'ha3:data=16'b1110111111111111;//STATE:24	SEG:3	COUNTER:163	
		10'ha4:data=16'b0010101010101011;//STATE:24	SEG:4	COUNTER:164	
		10'ha5:data=16'b1010101010001110;//STATE:24	SEG:5	COUNTER:165	
		10'ha6:data=16'b1011100011100011;//STATE:24	SEG:6	COUNTER:166	
		10'ha7:data=16'b1000000000000000;//STATE:24	SEG:7	COUNTER:167	
		10'ha8:data=16'b1001000010000001;//STATE:25	SEG:1	COUNTER:168	
		10'ha9:data=16'b0000000011111111;//STATE:25	SEG:2	COUNTER:169	
		10'haa:data=16'b1110111111111111;//STATE:25	SEG:3	COUNTER:170	
		10'hab:data=16'b0110101010101011;//STATE:25	SEG:4	COUNTER:171	
		10'hac:data=16'b1010101010101110;//STATE:25	SEG:5	COUNTER:172	
		10'had:data=16'b1011100011100011;//STATE:25	SEG:6	COUNTER:173	
		10'hae:data=16'b1001000000000000;//STATE:25	SEG:7	COUNTER:174	
		10'haf:data=16'b1001000010000001;//STATE:26	SEG:1	COUNTER:175	
		10'hb0:data=16'b0000000010111111;//STATE:26	SEG:2	COUNTER:176	
		10'hb1:data=16'b1110111111111111;//STATE:26	SEG:3	COUNTER:177	
		10'hb2:data=16'b0111101010101011;//STATE:26	SEG:4	COUNTER:178	
		10'hb3:data=16'b1010101010101010;//STATE:26	SEG:5	COUNTER:179	
		10'hb4:data=16'b1011100011100011;//STATE:26	SEG:6	COUNTER:180	
		10'hb5:data=16'b1001000000000000;//STATE:26	SEG:7	COUNTER:181	
		10'hb6:data=16'b1001000010000001;//STATE:27	SEG:1	COUNTER:182	
		10'hb7:data=16'b0000000010011111;//STATE:27	SEG:2	COUNTER:183	
		10'hb8:data=16'b1110111111111111;//STATE:27	SEG:3	COUNTER:184	
		10'hb9:data=16'b0111111010101011;//STATE:27	SEG:4	COUNTER:185	
		10'hba:data=16'b1010101010101010;//STATE:27	SEG:5	COUNTER:186	
		10'hbb:data=16'b0011100011100011;//STATE:27	SEG:6	COUNTER:187	
		10'hbc:data=16'b1001000000000000;//STATE:27	SEG:7	COUNTER:188	
		10'hbd:data=16'b1001000010000001;//STATE:28	SEG:1	COUNTER:189	
		10'hbe:data=16'b0000000010001111;//STATE:28	SEG:2	COUNTER:190	
		10'hbf:data=16'b1110111111111111;//STATE:28	SEG:3	COUNTER:191	
		10'hc0:data=16'b0111111110101011;//STATE:28	SEG:4	COUNTER:192	
		10'hc1:data=16'b1010101010101010;//STATE:28	SEG:5	COUNTER:193	
		10'hc2:data=16'b0010100011100011;//STATE:28	SEG:6	COUNTER:194	
		10'hc3:data=16'b1001000000000000;//STATE:28	SEG:7	COUNTER:195	
		10'hc4:data=16'b1001000010000001;//STATE:29	SEG:1	COUNTER:196	
		10'hc5:data=16'b0000000010000111;//STATE:29	SEG:2	COUNTER:197	
		10'hc6:data=16'b1110111111111111;//STATE:29	SEG:3	COUNTER:198	
		10'hc7:data=16'b0111111111101011;//STATE:29	SEG:4	COUNTER:199	
		10'hc8:data=16'b1010101010101010;//STATE:29	SEG:5	COUNTER:200	
		10'hc9:data=16'b0010101011100011;//STATE:29	SEG:6	COUNTER:201	
		10'hca:data=16'b1001000000000000;//STATE:29	SEG:7	COUNTER:202	
		10'hcb:data=16'b1001000010000001;//STATE:30	SEG:1	COUNTER:203	
		10'hcc:data=16'b0000000010000011;//STATE:30	SEG:2	COUNTER:204	
		10'hcd:data=16'b1110111111111111;//STATE:30	SEG:3	COUNTER:205	
		10'hce:data=16'b0111111111111011;//STATE:30	SEG:4	COUNTER:206	
		10'hcf:data=16'b1010101010101010;//STATE:30	SEG:5	COUNTER:207	
		10'hd0:data=16'b0010101010100011;//STATE:30	SEG:6	COUNTER:208	
		10'hd1:data=16'b1001000000000000;//STATE:30	SEG:7	COUNTER:209	
		10'hd2:data=16'b1001000010000001;//STATE:31	SEG:1	COUNTER:210	
		10'hd3:data=16'b0000000010000001;//STATE:31	SEG:2	COUNTER:211	
		10'hd4:data=16'b1110111111111111;//STATE:31	SEG:3	COUNTER:212	
		10'hd5:data=16'b0111111111111111;//STATE:31	SEG:4	COUNTER:213	
		10'hd6:data=16'b1010101010101010;//STATE:31	SEG:5	COUNTER:214	
		10'hd7:data=16'b0010101010101011;//STATE:31	SEG:6	COUNTER:215	
		10'hd8:data=16'b1001000000000000;//STATE:31	SEG:7	COUNTER:216	
		10'hd9:data=16'b1001000010000001;//STATE:32	SEG:1	COUNTER:217	
		10'hda:data=16'b0000000010000000;//STATE:32	SEG:2	COUNTER:218	
		10'hdb:data=16'b1110111111111111;//STATE:32	SEG:3	COUNTER:219	
		10'hdc:data=16'b0111111111111110;//STATE:32	SEG:4	COUNTER:220	
		10'hdd:data=16'b1010101010101010;//STATE:32	SEG:5	COUNTER:221	
		10'hde:data=16'b0010101010101010;//STATE:32	SEG:6	COUNTER:222	
		10'hdf:data=16'b1001000000000000;//STATE:32	SEG:7	COUNTER:223	
		10'he0:data=16'b1001000010000001;//STATE:33	SEG:1	COUNTER:224	
		10'he1:data=16'b0000000010000000;//STATE:33	SEG:2	COUNTER:225	
		10'he2:data=16'b0110111111111111;//STATE:33	SEG:3	COUNTER:226	
		10'he3:data=16'b0111111111111110;//STATE:33	SEG:4	COUNTER:227	
		10'he4:data=16'b1110101010101010;//STATE:33	SEG:5	COUNTER:228	
		10'he5:data=16'b0010101010101010;//STATE:33	SEG:6	COUNTER:229	
		10'he6:data=16'b1011000000000000;//STATE:33	SEG:7	COUNTER:230	
		10'he7:data=16'b1001000010000001;//STATE:34	SEG:1	COUNTER:231	
		10'he8:data=16'b0000000010000000;//STATE:34	SEG:2	COUNTER:232	
		10'he9:data=16'b0010111111111111;//STATE:34	SEG:3	COUNTER:233	
		10'hea:data=16'b0111111111111110;//STATE:34	SEG:4	COUNTER:234	
		10'heb:data=16'b1111101010101010;//STATE:34	SEG:5	COUNTER:235	
		10'hec:data=16'b0010101010101010;//STATE:34	SEG:6	COUNTER:236	
		10'hed:data=16'b1011000000000000;//STATE:34	SEG:7	COUNTER:237	
		10'hee:data=16'b1001000010000001;//STATE:35	SEG:1	COUNTER:238	
		10'hef:data=16'b0000000010000000;//STATE:35	SEG:2	COUNTER:239	
		10'hf0:data=16'b0000111111111111;//STATE:35	SEG:3	COUNTER:240	
		10'hf1:data=16'b0111111111111110;//STATE:35	SEG:4	COUNTER:241	
		10'hf2:data=16'b1111111010101010;//STATE:35	SEG:5	COUNTER:242	
		10'hf3:data=16'b0010101010101010;//STATE:35	SEG:6	COUNTER:243	
		10'hf4:data=16'b1011000000000000;//STATE:35	SEG:7	COUNTER:244	
		10'hf5:data=16'b1001000010000001;//STATE:36	SEG:1	COUNTER:245	
		10'hf6:data=16'b0000000010000000;//STATE:36	SEG:2	COUNTER:246	
		10'hf7:data=16'b0001111111111111;//STATE:36	SEG:3	COUNTER:247	
		10'hf8:data=16'b0111111111111110;//STATE:36	SEG:4	COUNTER:248	
		10'hf9:data=16'b1111111110101010;//STATE:36	SEG:5	COUNTER:249	
		10'hfa:data=16'b0010101010101010;//STATE:36	SEG:6	COUNTER:250	
		10'hfb:data=16'b1011000000000000;//STATE:36	SEG:7	COUNTER:251	
		10'hfc:data=16'b1001000010000001;//STATE:37	SEG:1	COUNTER:252	
		10'hfd:data=16'b0000000010000000;//STATE:37	SEG:2	COUNTER:253	
		10'hfe:data=16'b0001011111111111;//STATE:37	SEG:3	COUNTER:254	
		10'hff:data=16'b0111111111111110;//STATE:37	SEG:4	COUNTER:255	
		10'h100:data=16'b1111111111101010;//STATE:37	SEG:5	COUNTER:256	
		10'h101:data=16'b0010101010101010;//STATE:37	SEG:6	COUNTER:257	
		10'h102:data=16'b1011000000000000;//STATE:37	SEG:7	COUNTER:258	
		10'h103:data=16'b1001000010000001;//STATE:38	SEG:1	COUNTER:259	
		10'h104:data=16'b0000000010000000;//STATE:38	SEG:2	COUNTER:260	
		10'h105:data=16'b0001001111111111;//STATE:38	SEG:3	COUNTER:261	
		10'h106:data=16'b0111111111111110;//STATE:38	SEG:4	COUNTER:262	
		10'h107:data=16'b1111111111111010;//STATE:38	SEG:5	COUNTER:263	
		10'h108:data=16'b0010101010101010;//STATE:38	SEG:6	COUNTER:264	
		10'h109:data=16'b1011000000000000;//STATE:38	SEG:7	COUNTER:265	
		10'h10a:data=16'b1001000010000001;//STATE:39	SEG:1	COUNTER:266	
		10'h10b:data=16'b0000000010000000;//STATE:39	SEG:2	COUNTER:267	
		10'h10c:data=16'b0001000111111111;//STATE:39	SEG:3	COUNTER:268	
		10'h10d:data=16'b0111111111111110;//STATE:39	SEG:4	COUNTER:269	
		10'h10e:data=16'b1111111111111110;//STATE:39	SEG:5	COUNTER:270	
		10'h10f:data=16'b0010101010101010;//STATE:39	SEG:6	COUNTER:271	
		10'h110:data=16'b1011000000000000;//STATE:39	SEG:7	COUNTER:272	
		10'h111:data=16'b1001000010000001;//STATE:40	SEG:1	COUNTER:273	
		10'h112:data=16'b0000000010000000;//STATE:40	SEG:2	COUNTER:274	
		10'h113:data=16'b0001000011111111;//STATE:40	SEG:3	COUNTER:275	
		10'h114:data=16'b0111111111111110;//STATE:40	SEG:4	COUNTER:276	
		10'h115:data=16'b1111111111111111;//STATE:40	SEG:5	COUNTER:277	
		10'h116:data=16'b0010101010101010;//STATE:40	SEG:6	COUNTER:278	
		10'h117:data=16'b1011000000000000;//STATE:40	SEG:7	COUNTER:279	
		10'h118:data=16'b1001000010000001;//STATE:41	SEG:1	COUNTER:280	
		10'h119:data=16'b0000000010000000;//STATE:41	SEG:2	COUNTER:281	
		10'h11a:data=16'b0001000001111111;//STATE:41	SEG:3	COUNTER:282	
		10'h11b:data=16'b0111111111111110;//STATE:41	SEG:4	COUNTER:283	
		10'h11c:data=16'b1111111111111111;//STATE:41	SEG:5	COUNTER:284	
		10'h11d:data=16'b0110101010101010;//STATE:41	SEG:6	COUNTER:285	
		10'h11e:data=16'b1011000000000000;//STATE:41	SEG:7	COUNTER:286	
		10'h11f:data=16'b1001000010000001;//STATE:42	SEG:1	COUNTER:287	
		10'h120:data=16'b0000000010000000;//STATE:42	SEG:2	COUNTER:288	
		10'h121:data=16'b0001000000111111;//STATE:42	SEG:3	COUNTER:289	
		10'h122:data=16'b0111111111111110;//STATE:42	SEG:4	COUNTER:290	
		10'h123:data=16'b1111111111111111;//STATE:42	SEG:5	COUNTER:291	
		10'h124:data=16'b0111101010101010;//STATE:42	SEG:6	COUNTER:292	
		10'h125:data=16'b1011000000000000;//STATE:42	SEG:7	COUNTER:293	
		10'h126:data=16'b1001000010000001;//STATE:43	SEG:1	COUNTER:294	
		10'h127:data=16'b0000000010000000;//STATE:43	SEG:2	COUNTER:295	
		10'h128:data=16'b0001000000011111;//STATE:43	SEG:3	COUNTER:296	
		10'h129:data=16'b0111111111111110;//STATE:43	SEG:4	COUNTER:297	
		10'h12a:data=16'b1111111111111111;//STATE:43	SEG:5	COUNTER:298	
		10'h12b:data=16'b0111111010101010;//STATE:43	SEG:6	COUNTER:299	
		10'h12c:data=16'b1011000000000000;//STATE:43	SEG:7	COUNTER:300	
		10'h12d:data=16'b1001000010000001;//STATE:44	SEG:1	COUNTER:301	
		10'h12e:data=16'b0000000010000000;//STATE:44	SEG:2	COUNTER:302	
		10'h12f:data=16'b0001000000001111;//STATE:44	SEG:3	COUNTER:303	
		10'h130:data=16'b0111111111111110;//STATE:44	SEG:4	COUNTER:304	
		10'h131:data=16'b1111111111111111;//STATE:44	SEG:5	COUNTER:305	
		10'h132:data=16'b0111111110101010;//STATE:44	SEG:6	COUNTER:306	
		10'h133:data=16'b1011000000000000;//STATE:44	SEG:7	COUNTER:307	
		10'h134:data=16'b1001000010000001;//STATE:45	SEG:1	COUNTER:308	
		10'h135:data=16'b0000000010000000;//STATE:45	SEG:2	COUNTER:309	
		10'h136:data=16'b0001000000000111;//STATE:45	SEG:3	COUNTER:310	
		10'h137:data=16'b0111111111111110;//STATE:45	SEG:4	COUNTER:311	
		10'h138:data=16'b1111111111111111;//STATE:45	SEG:5	COUNTER:312	
		10'h139:data=16'b0111111111101010;//STATE:45	SEG:6	COUNTER:313	
		10'h13a:data=16'b1011000000000000;//STATE:45	SEG:7	COUNTER:314	
		10'h13b:data=16'b1001000010000001;//STATE:46	SEG:1	COUNTER:315	
		10'h13c:data=16'b0000000010000000;//STATE:46	SEG:2	COUNTER:316	
		10'h13d:data=16'b0001000000000011;//STATE:46	SEG:3	COUNTER:317	
		10'h13e:data=16'b0111111111111110;//STATE:46	SEG:4	COUNTER:318	
		10'h13f:data=16'b1111111111111111;//STATE:46	SEG:5	COUNTER:319	
		10'h140:data=16'b0111111111111010;//STATE:46	SEG:6	COUNTER:320	
		10'h141:data=16'b1011000000000000;//STATE:46	SEG:7	COUNTER:321	
		10'h142:data=16'b1001000010000001;//STATE:47	SEG:1	COUNTER:322	
		10'h143:data=16'b0000000010000000;//STATE:47	SEG:2	COUNTER:323	
		10'h144:data=16'b0001000000000001;//STATE:47	SEG:3	COUNTER:324	
		10'h145:data=16'b0111111111111110;//STATE:47	SEG:4	COUNTER:325	
		10'h146:data=16'b1111111111111111;//STATE:47	SEG:5	COUNTER:326	
		10'h147:data=16'b0111111111111110;//STATE:47	SEG:6	COUNTER:327	
		10'h148:data=16'b1011000000000000;//STATE:47	SEG:7	COUNTER:328	
		10'h149:data=16'b1001000010000001;//STATE:48	SEG:1	COUNTER:329	
		10'h14a:data=16'b0000000010000000;//STATE:48	SEG:2	COUNTER:330	
		10'h14b:data=16'b0001000000000000;//STATE:48	SEG:3	COUNTER:331	
		10'h14c:data=16'b0111111111111110;//STATE:48	SEG:4	COUNTER:332	
		10'h14d:data=16'b1111111111111111;//STATE:48	SEG:5	COUNTER:333	
		10'h14e:data=16'b0111111111111111;//STATE:48	SEG:6	COUNTER:334	
		10'h14f:data=16'b1011000000000000;//STATE:48	SEG:7	COUNTER:335	
		10'h150:data=16'b1001000010000001;//STATE:49	SEG:1	COUNTER:336	
		10'h151:data=16'b0000000010000000;//STATE:49	SEG:2	COUNTER:337	
		10'h152:data=16'b0001000000000000;//STATE:49	SEG:3	COUNTER:338	
		10'h153:data=16'b1111111111111110;//STATE:49	SEG:4	COUNTER:339	
		10'h154:data=16'b1111111111111111;//STATE:49	SEG:5	COUNTER:340	
		10'h155:data=16'b0111111111111111;//STATE:49	SEG:6	COUNTER:341	
		10'h156:data=16'b1111000000000000;//STATE:49	SEG:7	COUNTER:342	
		10'h157:data=16'b1001000010000001;//STATE:50	SEG:1	COUNTER:343	
		10'h158:data=16'b0000000010000000;//STATE:50	SEG:2	COUNTER:344	
		10'h159:data=16'b0001000000000000;//STATE:50	SEG:3	COUNTER:345	
		10'h15a:data=16'b1011111111111110;//STATE:50	SEG:4	COUNTER:346	
		10'h15b:data=16'b1111111111111111;//STATE:50	SEG:5	COUNTER:347	
		10'h15c:data=16'b0111111111111111;//STATE:50	SEG:6	COUNTER:348	
		10'h15d:data=16'b1110000000000000;//STATE:50	SEG:7	COUNTER:349	
		10'h15e:data=16'b1001000010000001;//STATE:51	SEG:1	COUNTER:350	
		10'h15f:data=16'b0000000010000000;//STATE:51	SEG:2	COUNTER:351	
		10'h160:data=16'b0001000000000000;//STATE:51	SEG:3	COUNTER:352	
		10'h161:data=16'b1001111111111110;//STATE:51	SEG:4	COUNTER:353	
		10'h162:data=16'b1111111111111111;//STATE:51	SEG:5	COUNTER:354	
		10'h163:data=16'b0111111111111111;//STATE:51	SEG:6	COUNTER:355	
		10'h164:data=16'b1110000000000000;//STATE:51	SEG:7	COUNTER:356	
		10'h165:data=16'b1001000010000001;//STATE:52	SEG:1	COUNTER:357	
		10'h166:data=16'b0000000010000000;//STATE:52	SEG:2	COUNTER:358	
		10'h167:data=16'b0001000000000000;//STATE:52	SEG:3	COUNTER:359	
		10'h168:data=16'b1000111111111110;//STATE:52	SEG:4	COUNTER:360	
		10'h169:data=16'b1111111111111111;//STATE:52	SEG:5	COUNTER:361	
		10'h16a:data=16'b0111111111111111;//STATE:52	SEG:6	COUNTER:362	
		10'h16b:data=16'b1110000000000000;//STATE:52	SEG:7	COUNTER:363	
		10'h16c:data=16'b1001000010000001;//STATE:53	SEG:1	COUNTER:364	
		10'h16d:data=16'b0000000010000000;//STATE:53	SEG:2	COUNTER:365	
		10'h16e:data=16'b0001000000000000;//STATE:53	SEG:3	COUNTER:366	
		10'h16f:data=16'b1000011111111110;//STATE:53	SEG:4	COUNTER:367	
		10'h170:data=16'b1111111111111111;//STATE:53	SEG:5	COUNTER:368	
		10'h171:data=16'b0111111111111111;//STATE:53	SEG:6	COUNTER:369	
		10'h172:data=16'b1110000000000000;//STATE:53	SEG:7	COUNTER:370	
		10'h173:data=16'b1001000010000001;//STATE:54	SEG:1	COUNTER:371	
		10'h174:data=16'b0000000010000000;//STATE:54	SEG:2	COUNTER:372	
		10'h175:data=16'b0001000000000000;//STATE:54	SEG:3	COUNTER:373	
		10'h176:data=16'b1000001111111110;//STATE:54	SEG:4	COUNTER:374	
		10'h177:data=16'b1111111111111111;//STATE:54	SEG:5	COUNTER:375	
		10'h178:data=16'b0111111111111111;//STATE:54	SEG:6	COUNTER:376	
		10'h179:data=16'b1110000000000000;//STATE:54	SEG:7	COUNTER:377	
		10'h17a:data=16'b1001000010000001;//STATE:55	SEG:1	COUNTER:378	
		10'h17b:data=16'b0000000010000000;//STATE:55	SEG:2	COUNTER:379	
		10'h17c:data=16'b0001000000000000;//STATE:55	SEG:3	COUNTER:380	
		10'h17d:data=16'b1000000111111110;//STATE:55	SEG:4	COUNTER:381	
		10'h17e:data=16'b1111111111111111;//STATE:55	SEG:5	COUNTER:382	
		10'h17f:data=16'b0111111111111111;//STATE:55	SEG:6	COUNTER:383	
		10'h180:data=16'b1110000000000000;//STATE:55	SEG:7	COUNTER:384	
		10'h181:data=16'b1001000010000001;//STATE:56	SEG:1	COUNTER:385	
		10'h182:data=16'b0000000010000000;//STATE:56	SEG:2	COUNTER:386	
		10'h183:data=16'b0001000000000000;//STATE:56	SEG:3	COUNTER:387	
		10'h184:data=16'b1000000011111110;//STATE:56	SEG:4	COUNTER:388	
		10'h185:data=16'b1111111111111111;//STATE:56	SEG:5	COUNTER:389	
		10'h186:data=16'b0111111111111111;//STATE:56	SEG:6	COUNTER:390	
		10'h187:data=16'b1110000000000000;//STATE:56	SEG:7	COUNTER:391	
		10'h188:data=16'b1001000010000001;//STATE:57	SEG:1	COUNTER:392	
		10'h189:data=16'b0000000010000000;//STATE:57	SEG:2	COUNTER:393	
		10'h18a:data=16'b0001000000000000;//STATE:57	SEG:3	COUNTER:394	
		10'h18b:data=16'b1000000001111110;//STATE:57	SEG:4	COUNTER:395	
		10'h18c:data=16'b1111111111111111;//STATE:57	SEG:5	COUNTER:396	
		10'h18d:data=16'b0111111111111111;//STATE:57	SEG:6	COUNTER:397	
		10'h18e:data=16'b1110000000000000;//STATE:57	SEG:7	COUNTER:398	
		10'h18f:data=16'b1001000010000001;//STATE:58	SEG:1	COUNTER:399	
		10'h190:data=16'b0000000010000000;//STATE:58	SEG:2	COUNTER:400	
		10'h191:data=16'b0001000000000000;//STATE:58	SEG:3	COUNTER:401	
		10'h192:data=16'b1000000000111110;//STATE:58	SEG:4	COUNTER:402	
		10'h193:data=16'b1111111111111111;//STATE:58	SEG:5	COUNTER:403	
		10'h194:data=16'b0111111111111111;//STATE:58	SEG:6	COUNTER:404	
		10'h195:data=16'b1110000000000000;//STATE:58	SEG:7	COUNTER:405	
		10'h196:data=16'b1001000010000001;//STATE:59	SEG:1	COUNTER:406	
		10'h197:data=16'b0000000010000000;//STATE:59	SEG:2	COUNTER:407	
		10'h198:data=16'b0001000000000000;//STATE:59	SEG:3	COUNTER:408	
		10'h199:data=16'b1000000000011110;//STATE:59	SEG:4	COUNTER:409	
		10'h19a:data=16'b1111111111111111;//STATE:59	SEG:5	COUNTER:410	
		10'h19b:data=16'b0111111111111111;//STATE:59	SEG:6	COUNTER:411	
		10'h19c:data=16'b1110000000000000;//STATE:59	SEG:7	COUNTER:412	
		10'h19d:data=16'b1001000010000001;//STATE:60	SEG:1	COUNTER:413	
		10'h19e:data=16'b0000000010000000;//STATE:60	SEG:2	COUNTER:414	
		10'h19f:data=16'b0001000000000000;//STATE:60	SEG:3	COUNTER:415	
		10'h1a0:data=16'b1000000000001110;//STATE:60	SEG:4	COUNTER:416	
		10'h1a1:data=16'b1111111111111111;//STATE:60	SEG:5	COUNTER:417	
		10'h1a2:data=16'b0111111111111111;//STATE:60	SEG:6	COUNTER:418	
		10'h1a3:data=16'b1110000000000000;//STATE:60	SEG:7	COUNTER:419	
		10'h1a4:data=16'b1001000010000001;//STATE:61	SEG:1	COUNTER:420	
		10'h1a5:data=16'b0000000010000000;//STATE:61	SEG:2	COUNTER:421	
		10'h1a6:data=16'b0001000000000000;//STATE:61	SEG:3	COUNTER:422	
		10'h1a7:data=16'b1000000000000110;//STATE:61	SEG:4	COUNTER:423	
		10'h1a8:data=16'b1111111111111111;//STATE:61	SEG:5	COUNTER:424	
		10'h1a9:data=16'b0111111111111111;//STATE:61	SEG:6	COUNTER:425	
		10'h1aa:data=16'b1110000000000000;//STATE:61	SEG:7	COUNTER:426	
		10'h1ab:data=16'b1001000010000001;//STATE:62	SEG:1	COUNTER:427	
		10'h1ac:data=16'b0000000010000000;//STATE:62	SEG:2	COUNTER:428	
		10'h1ad:data=16'b0001000000000000;//STATE:62	SEG:3	COUNTER:429	
		10'h1ae:data=16'b1000000000000010;//STATE:62	SEG:4	COUNTER:430	
		10'h1af:data=16'b1111111111111111;//STATE:62	SEG:5	COUNTER:431	
		10'h1b0:data=16'b0111111111111111;//STATE:62	SEG:6	COUNTER:432	
		10'h1b1:data=16'b1110000000000000;//STATE:62	SEG:7	COUNTER:433	
		10'h1b2:data=16'b1001000010000001;//STATE:63	SEG:1	COUNTER:434	
		10'h1b3:data=16'b0000000010000000;//STATE:63	SEG:2	COUNTER:435	
		10'h1b4:data=16'b0001000000000000;//STATE:63	SEG:3	COUNTER:436	
		10'h1b5:data=16'b1000000000000000;//STATE:63	SEG:4	COUNTER:437	
		10'h1b6:data=16'b1111111111111111;//STATE:63	SEG:5	COUNTER:438	
		10'h1b7:data=16'b0111111111111111;//STATE:63	SEG:6	COUNTER:439	
		10'h1b8:data=16'b1110000000000000;//STATE:63	SEG:7	COUNTER:440	
		10'h1b9:data=16'b1001000010000001;//STATE:64	SEG:1	COUNTER:441	
		10'h1ba:data=16'b0000000010000000;//STATE:64	SEG:2	COUNTER:442	
		10'h1bb:data=16'b0001000000000000;//STATE:64	SEG:3	COUNTER:443	
		10'h1bc:data=16'b1000000000000001;//STATE:64	SEG:4	COUNTER:444	
		10'h1bd:data=16'b1111111111111111;//STATE:64	SEG:5	COUNTER:445	
		10'h1be:data=16'b0111111111111111;//STATE:64	SEG:6	COUNTER:446	
		10'h1bf:data=16'b1110000000000000;//STATE:64	SEG:7	COUNTER:447	
		10'h1c0:data=16'b1001000010000001;//STATE:65	SEG:1	COUNTER:448	
		10'h1c1:data=16'b0000000010000000;//STATE:65	SEG:2	COUNTER:449	
		10'h1c2:data=16'b0001000000000000;//STATE:65	SEG:3	COUNTER:450	
		10'h1c3:data=16'b1000000000000001;//STATE:65	SEG:4	COUNTER:451	
		10'h1c4:data=16'b0111111111111111;//STATE:65	SEG:5	COUNTER:452	
		10'h1c5:data=16'b0111111111111111;//STATE:65	SEG:6	COUNTER:453	
		10'h1c6:data=16'b1110000000000000;//STATE:65	SEG:7	COUNTER:454	
		10'h1c7:data=16'b1001000010000001;//STATE:66	SEG:1	COUNTER:455	
		10'h1c8:data=16'b0000000010000000;//STATE:66	SEG:2	COUNTER:456	
		10'h1c9:data=16'b0001000000000000;//STATE:66	SEG:3	COUNTER:457	
		10'h1ca:data=16'b1000000000000001;//STATE:66	SEG:4	COUNTER:458	
		10'h1cb:data=16'b0011111111111111;//STATE:66	SEG:5	COUNTER:459	
		10'h1cc:data=16'b0111111111111111;//STATE:66	SEG:6	COUNTER:460	
		10'h1cd:data=16'b1110000000000000;//STATE:66	SEG:7	COUNTER:461	
		10'h1ce:data=16'b1001000010000001;//STATE:67	SEG:1	COUNTER:462	
		10'h1cf:data=16'b0000000010000000;//STATE:67	SEG:2	COUNTER:463	
		10'h1d0:data=16'b0001000000000000;//STATE:67	SEG:3	COUNTER:464	
		10'h1d1:data=16'b1000000000000001;//STATE:67	SEG:4	COUNTER:465	
		10'h1d2:data=16'b0001111111111111;//STATE:67	SEG:5	COUNTER:466	
		10'h1d3:data=16'b0111111111111111;//STATE:67	SEG:6	COUNTER:467	
		10'h1d4:data=16'b1110000000000000;//STATE:67	SEG:7	COUNTER:468	
		10'h1d5:data=16'b1001000010000001;//STATE:68	SEG:1	COUNTER:469	
		10'h1d6:data=16'b0000000010000000;//STATE:68	SEG:2	COUNTER:470	
		10'h1d7:data=16'b0001000000000000;//STATE:68	SEG:3	COUNTER:471	
		10'h1d8:data=16'b1000000000000001;//STATE:68	SEG:4	COUNTER:472	
		10'h1d9:data=16'b0000111111111111;//STATE:68	SEG:5	COUNTER:473	
		10'h1da:data=16'b0111111111111111;//STATE:68	SEG:6	COUNTER:474	
		10'h1db:data=16'b1110000000000000;//STATE:68	SEG:7	COUNTER:475	
		10'h1dc:data=16'b1001000010000001;//STATE:69	SEG:1	COUNTER:476	
		10'h1dd:data=16'b0000000010000000;//STATE:69	SEG:2	COUNTER:477	
		10'h1de:data=16'b0001000000000000;//STATE:69	SEG:3	COUNTER:478	
		10'h1df:data=16'b1000000000000001;//STATE:69	SEG:4	COUNTER:479	
		10'h1e0:data=16'b0000011111111111;//STATE:69	SEG:5	COUNTER:480	
		10'h1e1:data=16'b0111111111111111;//STATE:69	SEG:6	COUNTER:481	
		10'h1e2:data=16'b1110000000000000;//STATE:69	SEG:7	COUNTER:482	
		10'h1e3:data=16'b1001000010000001;//STATE:70	SEG:1	COUNTER:483	
		10'h1e4:data=16'b0000000010000000;//STATE:70	SEG:2	COUNTER:484	
		10'h1e5:data=16'b0001000000000000;//STATE:70	SEG:3	COUNTER:485	
		10'h1e6:data=16'b1000000000000001;//STATE:70	SEG:4	COUNTER:486	
		10'h1e7:data=16'b0000001111111111;//STATE:70	SEG:5	COUNTER:487	
		10'h1e8:data=16'b0111111111111111;//STATE:70	SEG:6	COUNTER:488	
		10'h1e9:data=16'b1110000000000000;//STATE:70	SEG:7	COUNTER:489	
		10'h1ea:data=16'b1001000010000001;//STATE:71	SEG:1	COUNTER:490	
		10'h1eb:data=16'b0000000010000000;//STATE:71	SEG:2	COUNTER:491	
		10'h1ec:data=16'b0001000000000000;//STATE:71	SEG:3	COUNTER:492	
		10'h1ed:data=16'b1000000000000001;//STATE:71	SEG:4	COUNTER:493	
		10'h1ee:data=16'b0000000111111111;//STATE:71	SEG:5	COUNTER:494	
		10'h1ef:data=16'b0111111111111111;//STATE:71	SEG:6	COUNTER:495	
		10'h1f0:data=16'b1110000000000000;//STATE:71	SEG:7	COUNTER:496	
		10'h1f1:data=16'b1001000010000001;//STATE:72	SEG:1	COUNTER:497	
		10'h1f2:data=16'b0000000010000000;//STATE:72	SEG:2	COUNTER:498	
		10'h1f3:data=16'b0001000000000000;//STATE:72	SEG:3	COUNTER:499	
		10'h1f4:data=16'b1000000000000001;//STATE:72	SEG:4	COUNTER:500	
		10'h1f5:data=16'b0000000011111111;//STATE:72	SEG:5	COUNTER:501	
		10'h1f6:data=16'b0111111111111111;//STATE:72	SEG:6	COUNTER:502	
		10'h1f7:data=16'b1110000000000000;//STATE:72	SEG:7	COUNTER:503	
		10'h1f8:data=16'b1001000010000001;//STATE:73	SEG:1	COUNTER:504	
		10'h1f9:data=16'b0000000010000000;//STATE:73	SEG:2	COUNTER:505	
		10'h1fa:data=16'b0001000000000000;//STATE:73	SEG:3	COUNTER:506	
		10'h1fb:data=16'b1000000000000001;//STATE:73	SEG:4	COUNTER:507	
		10'h1fc:data=16'b0000000001111111;//STATE:73	SEG:5	COUNTER:508	
		10'h1fd:data=16'b0111111111111111;//STATE:73	SEG:6	COUNTER:509	
		10'h1fe:data=16'b1110000000000000;//STATE:73	SEG:7	COUNTER:510	
		10'h1ff:data=16'b1001000010000001;//STATE:74	SEG:1	COUNTER:511	
		10'h200:data=16'b0000000010000000;//STATE:74	SEG:2	COUNTER:512	
		10'h201:data=16'b0001000000000000;//STATE:74	SEG:3	COUNTER:513	
		10'h202:data=16'b1000000000000001;//STATE:74	SEG:4	COUNTER:514	
		10'h203:data=16'b0000000000111111;//STATE:74	SEG:5	COUNTER:515	
		10'h204:data=16'b0111111111111111;//STATE:74	SEG:6	COUNTER:516	
		10'h205:data=16'b1110000000000000;//STATE:74	SEG:7	COUNTER:517	
		10'h206:data=16'b1001000010000001;//STATE:75	SEG:1	COUNTER:518	
		10'h207:data=16'b0000000010000000;//STATE:75	SEG:2	COUNTER:519	
		10'h208:data=16'b0001000000000000;//STATE:75	SEG:3	COUNTER:520	
		10'h209:data=16'b1000000000000001;//STATE:75	SEG:4	COUNTER:521	
		10'h20a:data=16'b0000000000011111;//STATE:75	SEG:5	COUNTER:522	
		10'h20b:data=16'b0111111111111111;//STATE:75	SEG:6	COUNTER:523	
		10'h20c:data=16'b1110000000000000;//STATE:75	SEG:7	COUNTER:524	
		10'h20d:data=16'b1001000010000001;//STATE:76	SEG:1	COUNTER:525	
		10'h20e:data=16'b0000000010000000;//STATE:76	SEG:2	COUNTER:526	
		10'h20f:data=16'b0001000000000000;//STATE:76	SEG:3	COUNTER:527	
		10'h210:data=16'b1000000000000001;//STATE:76	SEG:4	COUNTER:528	
		10'h211:data=16'b0000000000001111;//STATE:76	SEG:5	COUNTER:529	
		10'h212:data=16'b0111111111111111;//STATE:76	SEG:6	COUNTER:530	
		10'h213:data=16'b1110000000000000;//STATE:76	SEG:7	COUNTER:531	
		10'h214:data=16'b1001000010000001;//STATE:77	SEG:1	COUNTER:532	
		10'h215:data=16'b0000000010000000;//STATE:77	SEG:2	COUNTER:533	
		10'h216:data=16'b0001000000000000;//STATE:77	SEG:3	COUNTER:534	
		10'h217:data=16'b1000000000000001;//STATE:77	SEG:4	COUNTER:535	
		10'h218:data=16'b0000000000000111;//STATE:77	SEG:5	COUNTER:536	
		10'h219:data=16'b0111111111111111;//STATE:77	SEG:6	COUNTER:537	
		10'h21a:data=16'b1110000000000000;//STATE:77	SEG:7	COUNTER:538	
		10'h21b:data=16'b1001000010000001;//STATE:78	SEG:1	COUNTER:539	
		10'h21c:data=16'b0000000010000000;//STATE:78	SEG:2	COUNTER:540	
		10'h21d:data=16'b0001000000000000;//STATE:78	SEG:3	COUNTER:541	
		10'h21e:data=16'b1000000000000001;//STATE:78	SEG:4	COUNTER:542	
		10'h21f:data=16'b0000000000000011;//STATE:78	SEG:5	COUNTER:543	
		10'h220:data=16'b0111111111111111;//STATE:78	SEG:6	COUNTER:544	
		10'h221:data=16'b1110000000000000;//STATE:78	SEG:7	COUNTER:545	
		10'h222:data=16'b1001000010000001;//STATE:79	SEG:1	COUNTER:546	
		10'h223:data=16'b0000000010000000;//STATE:79	SEG:2	COUNTER:547	
		10'h224:data=16'b0001000000000000;//STATE:79	SEG:3	COUNTER:548	
		10'h225:data=16'b1000000000000001;//STATE:79	SEG:4	COUNTER:549	
		10'h226:data=16'b0000000000000001;//STATE:79	SEG:5	COUNTER:550	
		10'h227:data=16'b0111111111111111;//STATE:79	SEG:6	COUNTER:551	
		10'h228:data=16'b1110000000000000;//STATE:79	SEG:7	COUNTER:552	
		10'h229:data=16'b1001000010000001;//STATE:80	SEG:1	COUNTER:553	
		10'h22a:data=16'b0000000010000000;//STATE:80	SEG:2	COUNTER:554	
		10'h22b:data=16'b0001000000000000;//STATE:80	SEG:3	COUNTER:555	
		10'h22c:data=16'b1000000000000001;//STATE:80	SEG:4	COUNTER:556	
		10'h22d:data=16'b0000000000000000;//STATE:80	SEG:5	COUNTER:557	
		10'h22e:data=16'b0111111111111111;//STATE:80	SEG:6	COUNTER:558	
		10'h22f:data=16'b1110000000000000;//STATE:80	SEG:7	COUNTER:559	
		10'h230:data=16'b1001000010000001;//STATE:81	SEG:1	COUNTER:560	
		10'h231:data=16'b0000000010000000;//STATE:81	SEG:2	COUNTER:561	
		10'h232:data=16'b0001000000000000;//STATE:81	SEG:3	COUNTER:562	
		10'h233:data=16'b1000000000000001;//STATE:81	SEG:4	COUNTER:563	
		10'h234:data=16'b0000000000000000;//STATE:81	SEG:5	COUNTER:564	
		10'h235:data=16'b1111111111111111;//STATE:81	SEG:6	COUNTER:565	
		10'h236:data=16'b1110000000000000;//STATE:81	SEG:7	COUNTER:566	
		10'h237:data=16'b1001000010000001;//STATE:82	SEG:1	COUNTER:567	
		10'h238:data=16'b0000000010000000;//STATE:82	SEG:2	COUNTER:568	
		10'h239:data=16'b0001000000000000;//STATE:82	SEG:3	COUNTER:569	
		10'h23a:data=16'b1000000000000001;//STATE:82	SEG:4	COUNTER:570	
		10'h23b:data=16'b0000000000000000;//STATE:82	SEG:5	COUNTER:571	
		10'h23c:data=16'b1011111111111111;//STATE:82	SEG:6	COUNTER:572	
		10'h23d:data=16'b1110000000000000;//STATE:82	SEG:7	COUNTER:573	
		10'h23e:data=16'b1001000010000001;//STATE:83	SEG:1	COUNTER:574	
		10'h23f:data=16'b0000000010000000;//STATE:83	SEG:2	COUNTER:575	
		10'h240:data=16'b0001000000000000;//STATE:83	SEG:3	COUNTER:576	
		10'h241:data=16'b1000000000000001;//STATE:83	SEG:4	COUNTER:577	
		10'h242:data=16'b0000000000000000;//STATE:83	SEG:5	COUNTER:578	
		10'h243:data=16'b1001111111111111;//STATE:83	SEG:6	COUNTER:579	
		10'h244:data=16'b1110000000000000;//STATE:83	SEG:7	COUNTER:580	
		10'h245:data=16'b1001000010000001;//STATE:84	SEG:1	COUNTER:581	
		10'h246:data=16'b0000000010000000;//STATE:84	SEG:2	COUNTER:582	
		10'h247:data=16'b0001000000000000;//STATE:84	SEG:3	COUNTER:583	
		10'h248:data=16'b1000000000000001;//STATE:84	SEG:4	COUNTER:584	
		10'h249:data=16'b0000000000000000;//STATE:84	SEG:5	COUNTER:585	
		10'h24a:data=16'b1000111111111111;//STATE:84	SEG:6	COUNTER:586	
		10'h24b:data=16'b1110000000000000;//STATE:84	SEG:7	COUNTER:587	
		10'h24c:data=16'b1001000010000001;//STATE:85	SEG:1	COUNTER:588	
		10'h24d:data=16'b0000000010000000;//STATE:85	SEG:2	COUNTER:589	
		10'h24e:data=16'b0001000000000000;//STATE:85	SEG:3	COUNTER:590	
		10'h24f:data=16'b1000000000000001;//STATE:85	SEG:4	COUNTER:591	
		10'h250:data=16'b0000000000000000;//STATE:85	SEG:5	COUNTER:592	
		10'h251:data=16'b1000011111111111;//STATE:85	SEG:6	COUNTER:593	
		10'h252:data=16'b1110000000000000;//STATE:85	SEG:7	COUNTER:594	
		10'h253:data=16'b1001000010000001;//STATE:86	SEG:1	COUNTER:595	
		10'h254:data=16'b0000000010000000;//STATE:86	SEG:2	COUNTER:596	
		10'h255:data=16'b0001000000000000;//STATE:86	SEG:3	COUNTER:597	
		10'h256:data=16'b1000000000000001;//STATE:86	SEG:4	COUNTER:598	
		10'h257:data=16'b0000000000000000;//STATE:86	SEG:5	COUNTER:599	
		10'h258:data=16'b1000001111111111;//STATE:86	SEG:6	COUNTER:600	
		10'h259:data=16'b1110000000000000;//STATE:86	SEG:7	COUNTER:601	
		10'h25a:data=16'b1001000010000001;//STATE:87	SEG:1	COUNTER:602	
		10'h25b:data=16'b0000000010000000;//STATE:87	SEG:2	COUNTER:603	
		10'h25c:data=16'b0001000000000000;//STATE:87	SEG:3	COUNTER:604	
		10'h25d:data=16'b1000000000000001;//STATE:87	SEG:4	COUNTER:605	
		10'h25e:data=16'b0000000000000000;//STATE:87	SEG:5	COUNTER:606	
		10'h25f:data=16'b1000000111111111;//STATE:87	SEG:6	COUNTER:607	
		10'h260:data=16'b1110000000000000;//STATE:87	SEG:7	COUNTER:608	
		10'h261:data=16'b1001000010000001;//STATE:88	SEG:1	COUNTER:609	
		10'h262:data=16'b0000000010000000;//STATE:88	SEG:2	COUNTER:610	
		10'h263:data=16'b0001000000000000;//STATE:88	SEG:3	COUNTER:611	
		10'h264:data=16'b1000000000000001;//STATE:88	SEG:4	COUNTER:612	
		10'h265:data=16'b0000000000000000;//STATE:88	SEG:5	COUNTER:613	
		10'h266:data=16'b1000000011111111;//STATE:88	SEG:6	COUNTER:614	
		10'h267:data=16'b1110000000000000;//STATE:88	SEG:7	COUNTER:615	
		10'h268:data=16'b1001000010000001;//STATE:89	SEG:1	COUNTER:616	
		10'h269:data=16'b0000000010000000;//STATE:89	SEG:2	COUNTER:617	
		10'h26a:data=16'b0001000000000000;//STATE:89	SEG:3	COUNTER:618	
		10'h26b:data=16'b1000000000000001;//STATE:89	SEG:4	COUNTER:619	
		10'h26c:data=16'b0000000000000000;//STATE:89	SEG:5	COUNTER:620	
		10'h26d:data=16'b1000000001111111;//STATE:89	SEG:6	COUNTER:621	
		10'h26e:data=16'b1110000000000000;//STATE:89	SEG:7	COUNTER:622	
		10'h26f:data=16'b1001000010000001;//STATE:90	SEG:1	COUNTER:623	
		10'h270:data=16'b0000000010000000;//STATE:90	SEG:2	COUNTER:624	
		10'h271:data=16'b0001000000000000;//STATE:90	SEG:3	COUNTER:625	
		10'h272:data=16'b1000000000000001;//STATE:90	SEG:4	COUNTER:626	
		10'h273:data=16'b0000000000000000;//STATE:90	SEG:5	COUNTER:627	
		10'h274:data=16'b1000000000111111;//STATE:90	SEG:6	COUNTER:628	
		10'h275:data=16'b1110000000000000;//STATE:90	SEG:7	COUNTER:629	
		10'h276:data=16'b1001000010000001;//STATE:91	SEG:1	COUNTER:630	
		10'h277:data=16'b0000000010000000;//STATE:91	SEG:2	COUNTER:631	
		10'h278:data=16'b0001000000000000;//STATE:91	SEG:3	COUNTER:632	
		10'h279:data=16'b1000000000000001;//STATE:91	SEG:4	COUNTER:633	
		10'h27a:data=16'b0000000000000000;//STATE:91	SEG:5	COUNTER:634	
		10'h27b:data=16'b1000000000011111;//STATE:91	SEG:6	COUNTER:635	
		10'h27c:data=16'b1110000000000000;//STATE:91	SEG:7	COUNTER:636	
		10'h27d:data=16'b1001000010000001;//STATE:92	SEG:1	COUNTER:637	
		10'h27e:data=16'b0000000010000000;//STATE:92	SEG:2	COUNTER:638	
		10'h27f:data=16'b0001000000000000;//STATE:92	SEG:3	COUNTER:639	
		10'h280:data=16'b1000000000000001;//STATE:92	SEG:4	COUNTER:640	
		10'h281:data=16'b0000000000000000;//STATE:92	SEG:5	COUNTER:641	
		10'h282:data=16'b1000000000001111;//STATE:92	SEG:6	COUNTER:642	
		10'h283:data=16'b1110000000000000;//STATE:92	SEG:7	COUNTER:643	
		10'h284:data=16'b1001000010000001;//STATE:93	SEG:1	COUNTER:644	
		10'h285:data=16'b0000000010000000;//STATE:93	SEG:2	COUNTER:645	
		10'h286:data=16'b0001000000000000;//STATE:93	SEG:3	COUNTER:646	
		10'h287:data=16'b1000000000000001;//STATE:93	SEG:4	COUNTER:647	
		10'h288:data=16'b0000000000000000;//STATE:93	SEG:5	COUNTER:648	
		10'h289:data=16'b1000000000000111;//STATE:93	SEG:6	COUNTER:649	
		10'h28a:data=16'b1110000000000000;//STATE:93	SEG:7	COUNTER:650	
		10'h28b:data=16'b1001000010000001;//STATE:94	SEG:1	COUNTER:651	
		10'h28c:data=16'b0000000010000000;//STATE:94	SEG:2	COUNTER:652	
		10'h28d:data=16'b0001000000000000;//STATE:94	SEG:3	COUNTER:653	
		10'h28e:data=16'b1000000000000001;//STATE:94	SEG:4	COUNTER:654	
		10'h28f:data=16'b0000000000000000;//STATE:94	SEG:5	COUNTER:655	
		10'h290:data=16'b1000000000000011;//STATE:94	SEG:6	COUNTER:656	
		10'h291:data=16'b1110000000000000;//STATE:94	SEG:7	COUNTER:657	
		10'h292:data=16'b1001000010000001;//STATE:95	SEG:1	COUNTER:658	
		10'h293:data=16'b0000000010000000;//STATE:95	SEG:2	COUNTER:659	
		10'h294:data=16'b0001000000000000;//STATE:95	SEG:3	COUNTER:660	
		10'h295:data=16'b1000000000000001;//STATE:95	SEG:4	COUNTER:661	
		10'h296:data=16'b0000000000000000;//STATE:95	SEG:5	COUNTER:662	
		10'h297:data=16'b1000000000000001;//STATE:95	SEG:6	COUNTER:663	
		10'h298:data=16'b1110000000000000;//STATE:95	SEG:7	COUNTER:664	
		10'h299:data=16'b1001000010000001;//STATE:96	SEG:1	COUNTER:665	
		10'h29a:data=16'b0000000010000000;//STATE:96	SEG:2	COUNTER:666	
		10'h29b:data=16'b0001000000000000;//STATE:96	SEG:3	COUNTER:667	
		10'h29c:data=16'b1000000000000001;//STATE:96	SEG:4	COUNTER:668	
		10'h29d:data=16'b0000000000000000;//STATE:96	SEG:5	COUNTER:669	
		10'h29e:data=16'b1000000000000000;//STATE:96	SEG:6	COUNTER:670	
		10'h29f:data=16'b1110000000000000;//STATE:96	SEG:7	COUNTER:671	
		10'h2a0:data=16'b1001000010000001;//STATE:97	SEG:1	COUNTER:672	
		10'h2a1:data=16'b0000000010000000;//STATE:97	SEG:2	COUNTER:673	
		10'h2a2:data=16'b0001000000000000;//STATE:97	SEG:3	COUNTER:674	
		10'h2a3:data=16'b1000000000000001;//STATE:97	SEG:4	COUNTER:675	
		10'h2a4:data=16'b0000000000000000;//STATE:97	SEG:5	COUNTER:676	
		10'h2a5:data=16'b1000000000000000;//STATE:97	SEG:6	COUNTER:677	
		10'h2a6:data=16'b0110000000000000;//STATE:97	SEG:7	COUNTER:678	
		10'h2a7:data=16'b1001000010000001;//STATE:98	SEG:1	COUNTER:679	
		10'h2a8:data=16'b0000000010000000;//STATE:98	SEG:2	COUNTER:680	
		10'h2a9:data=16'b0001000000000000;//STATE:98	SEG:3	COUNTER:681	
		10'h2aa:data=16'b1000000000000001;//STATE:98	SEG:4	COUNTER:682	
		10'h2ab:data=16'b0000000000000000;//STATE:98	SEG:5	COUNTER:683	
		10'h2ac:data=16'b1000000000000000;//STATE:98	SEG:6	COUNTER:684	
		10'h2ad:data=16'b0010000000000000;//STATE:98	SEG:7	COUNTER:685	
		10'h2ae:data=16'b1001000010000001;//STATE:99	SEG:1	COUNTER:686	
		10'h2af:data=16'b0000000010000000;//STATE:99	SEG:2	COUNTER:687	
		10'h2b0:data=16'b0001000000000000;//STATE:99	SEG:3	COUNTER:688	
		10'h2b1:data=16'b1000000000000001;//STATE:99	SEG:4	COUNTER:689	
		10'h2b2:data=16'b0000000000000000;//STATE:99	SEG:5	COUNTER:690	
		10'h2b3:data=16'b1000000000000000;//STATE:99	SEG:6	COUNTER:691	
		10'h2b4:data=16'b0000000000000000;//STATE:99	SEG:7	COUNTER:692	
		10'h2b5:data=16'b1001000010000001;//STATE:100	SEG:1	COUNTER:693	
		10'h2b6:data=16'b0000000010000000;//STATE:100	SEG:2	COUNTER:694	
		10'h2b7:data=16'b0001000000000000;//STATE:100	SEG:3	COUNTER:695	
		10'h2b8:data=16'b1000000000000001;//STATE:100	SEG:4	COUNTER:696	
		10'h2b9:data=16'b0000000000000000;//STATE:100	SEG:5	COUNTER:697	
		10'h2ba:data=16'b1000000000000000;//STATE:100	SEG:6	COUNTER:698	
		10'h2bb:data=16'b0001000000000000;//STATE:100	SEG:7	COUNTER:699	
        default:data=0;
    endcase
end
endmodule
