
`timescale 1us/10ns
module BPartCounter(
    input trigger,
    input SysRst,
    output reg [9:0] address
);

wire U1Carry;
wire U2Carry;
wire ResetSignal;
wire [3:0]U1Q;
wire [3:0]U2Q;
wire [3:0]U3Q;

HC74160 U1(
    ._LD(1),
    ._RD(ResetSignal),
    .D(4'b0),
    .CLK(trigger),
    .EP(1),
    .ET(1),
    .Q(U1Q),
    .C(U1Carry)
);
HC74160 U2(
    ._LD(1),
    ._RD(ResetSignal),
    .D(4'b0),
    .CLK(U1Carry),
    .EP(1),
    .ET(1),
    .Q(U2Q),
    .C(U2Carry)
);
HC74160 U3(
    ._LD(1),
    ._RD(ResetSignal),
    .D(4'b0),
    .CLK(U2Carry),
    .EP(1),
    .ET(1),
    .Q(U3Q),
    .C(U3Carry)
); 
wire asyncClrSignal;
assign asyncClrSignal = ~&{((~U1Q[0])&(~U1Q[1])&(~U1Q[2])&(~U1Q[3])),((~U2Q[0])&(~U2Q[1])&(~U2Q[2])&(~U2Q[3])),(U3Q[0]&U3Q[1]&U3Q[2]&(~U3Q[3]))};
and#(2)(ResetSignal ,(~SysRst) , asyncClrSignal);

always @(*) begin
    case({U3Q,U2Q,U1Q})
        //
        //12'b00001
//for i in range(0,700):
//    st='%03d'%i
//    print("\t\t12'b{0:04b}{1:04b}{2:04b}:address=10'd{3:d};".format(int(st[0]),int(st[1]),int(st[2]),i))
		12'b000000000000:address=10'd0;
		12'b000000000001:address=10'd1;
		12'b000000000010:address=10'd2;
		12'b000000000011:address=10'd3;
		12'b000000000100:address=10'd4;
		12'b000000000101:address=10'd5;
		12'b000000000110:address=10'd6;
		12'b000000000111:address=10'd7;
		12'b000000001000:address=10'd8;
		12'b000000001001:address=10'd9;
		12'b000000010000:address=10'd10;
		12'b000000010001:address=10'd11;
		12'b000000010010:address=10'd12;
		12'b000000010011:address=10'd13;
		12'b000000010100:address=10'd14;
		12'b000000010101:address=10'd15;
		12'b000000010110:address=10'd16;
		12'b000000010111:address=10'd17;
		12'b000000011000:address=10'd18;
		12'b000000011001:address=10'd19;
		12'b000000100000:address=10'd20;
		12'b000000100001:address=10'd21;
		12'b000000100010:address=10'd22;
		12'b000000100011:address=10'd23;
		12'b000000100100:address=10'd24;
		12'b000000100101:address=10'd25;
		12'b000000100110:address=10'd26;
		12'b000000100111:address=10'd27;
		12'b000000101000:address=10'd28;
		12'b000000101001:address=10'd29;
		12'b000000110000:address=10'd30;
		12'b000000110001:address=10'd31;
		12'b000000110010:address=10'd32;
		12'b000000110011:address=10'd33;
		12'b000000110100:address=10'd34;
		12'b000000110101:address=10'd35;
		12'b000000110110:address=10'd36;
		12'b000000110111:address=10'd37;
		12'b000000111000:address=10'd38;
		12'b000000111001:address=10'd39;
		12'b000001000000:address=10'd40;
		12'b000001000001:address=10'd41;
		12'b000001000010:address=10'd42;
		12'b000001000011:address=10'd43;
		12'b000001000100:address=10'd44;
		12'b000001000101:address=10'd45;
		12'b000001000110:address=10'd46;
		12'b000001000111:address=10'd47;
		12'b000001001000:address=10'd48;
		12'b000001001001:address=10'd49;
		12'b000001010000:address=10'd50;
		12'b000001010001:address=10'd51;
		12'b000001010010:address=10'd52;
		12'b000001010011:address=10'd53;
		12'b000001010100:address=10'd54;
		12'b000001010101:address=10'd55;
		12'b000001010110:address=10'd56;
		12'b000001010111:address=10'd57;
		12'b000001011000:address=10'd58;
		12'b000001011001:address=10'd59;
		12'b000001100000:address=10'd60;
		12'b000001100001:address=10'd61;
		12'b000001100010:address=10'd62;
		12'b000001100011:address=10'd63;
		12'b000001100100:address=10'd64;
		12'b000001100101:address=10'd65;
		12'b000001100110:address=10'd66;
		12'b000001100111:address=10'd67;
		12'b000001101000:address=10'd68;
		12'b000001101001:address=10'd69;
		12'b000001110000:address=10'd70;
		12'b000001110001:address=10'd71;
		12'b000001110010:address=10'd72;
		12'b000001110011:address=10'd73;
		12'b000001110100:address=10'd74;
		12'b000001110101:address=10'd75;
		12'b000001110110:address=10'd76;
		12'b000001110111:address=10'd77;
		12'b000001111000:address=10'd78;
		12'b000001111001:address=10'd79;
		12'b000010000000:address=10'd80;
		12'b000010000001:address=10'd81;
		12'b000010000010:address=10'd82;
		12'b000010000011:address=10'd83;
		12'b000010000100:address=10'd84;
		12'b000010000101:address=10'd85;
		12'b000010000110:address=10'd86;
		12'b000010000111:address=10'd87;
		12'b000010001000:address=10'd88;
		12'b000010001001:address=10'd89;
		12'b000010010000:address=10'd90;
		12'b000010010001:address=10'd91;
		12'b000010010010:address=10'd92;
		12'b000010010011:address=10'd93;
		12'b000010010100:address=10'd94;
		12'b000010010101:address=10'd95;
		12'b000010010110:address=10'd96;
		12'b000010010111:address=10'd97;
		12'b000010011000:address=10'd98;
		12'b000010011001:address=10'd99;
		12'b000100000000:address=10'd100;
		12'b000100000001:address=10'd101;
		12'b000100000010:address=10'd102;
		12'b000100000011:address=10'd103;
		12'b000100000100:address=10'd104;
		12'b000100000101:address=10'd105;
		12'b000100000110:address=10'd106;
		12'b000100000111:address=10'd107;
		12'b000100001000:address=10'd108;
		12'b000100001001:address=10'd109;
		12'b000100010000:address=10'd110;
		12'b000100010001:address=10'd111;
		12'b000100010010:address=10'd112;
		12'b000100010011:address=10'd113;
		12'b000100010100:address=10'd114;
		12'b000100010101:address=10'd115;
		12'b000100010110:address=10'd116;
		12'b000100010111:address=10'd117;
		12'b000100011000:address=10'd118;
		12'b000100011001:address=10'd119;
		12'b000100100000:address=10'd120;
		12'b000100100001:address=10'd121;
		12'b000100100010:address=10'd122;
		12'b000100100011:address=10'd123;
		12'b000100100100:address=10'd124;
		12'b000100100101:address=10'd125;
		12'b000100100110:address=10'd126;
		12'b000100100111:address=10'd127;
		12'b000100101000:address=10'd128;
		12'b000100101001:address=10'd129;
		12'b000100110000:address=10'd130;
		12'b000100110001:address=10'd131;
		12'b000100110010:address=10'd132;
		12'b000100110011:address=10'd133;
		12'b000100110100:address=10'd134;
		12'b000100110101:address=10'd135;
		12'b000100110110:address=10'd136;
		12'b000100110111:address=10'd137;
		12'b000100111000:address=10'd138;
		12'b000100111001:address=10'd139;
		12'b000101000000:address=10'd140;
		12'b000101000001:address=10'd141;
		12'b000101000010:address=10'd142;
		12'b000101000011:address=10'd143;
		12'b000101000100:address=10'd144;
		12'b000101000101:address=10'd145;
		12'b000101000110:address=10'd146;
		12'b000101000111:address=10'd147;
		12'b000101001000:address=10'd148;
		12'b000101001001:address=10'd149;
		12'b000101010000:address=10'd150;
		12'b000101010001:address=10'd151;
		12'b000101010010:address=10'd152;
		12'b000101010011:address=10'd153;
		12'b000101010100:address=10'd154;
		12'b000101010101:address=10'd155;
		12'b000101010110:address=10'd156;
		12'b000101010111:address=10'd157;
		12'b000101011000:address=10'd158;
		12'b000101011001:address=10'd159;
		12'b000101100000:address=10'd160;
		12'b000101100001:address=10'd161;
		12'b000101100010:address=10'd162;
		12'b000101100011:address=10'd163;
		12'b000101100100:address=10'd164;
		12'b000101100101:address=10'd165;
		12'b000101100110:address=10'd166;
		12'b000101100111:address=10'd167;
		12'b000101101000:address=10'd168;
		12'b000101101001:address=10'd169;
		12'b000101110000:address=10'd170;
		12'b000101110001:address=10'd171;
		12'b000101110010:address=10'd172;
		12'b000101110011:address=10'd173;
		12'b000101110100:address=10'd174;
		12'b000101110101:address=10'd175;
		12'b000101110110:address=10'd176;
		12'b000101110111:address=10'd177;
		12'b000101111000:address=10'd178;
		12'b000101111001:address=10'd179;
		12'b000110000000:address=10'd180;
		12'b000110000001:address=10'd181;
		12'b000110000010:address=10'd182;
		12'b000110000011:address=10'd183;
		12'b000110000100:address=10'd184;
		12'b000110000101:address=10'd185;
		12'b000110000110:address=10'd186;
		12'b000110000111:address=10'd187;
		12'b000110001000:address=10'd188;
		12'b000110001001:address=10'd189;
		12'b000110010000:address=10'd190;
		12'b000110010001:address=10'd191;
		12'b000110010010:address=10'd192;
		12'b000110010011:address=10'd193;
		12'b000110010100:address=10'd194;
		12'b000110010101:address=10'd195;
		12'b000110010110:address=10'd196;
		12'b000110010111:address=10'd197;
		12'b000110011000:address=10'd198;
		12'b000110011001:address=10'd199;
		12'b001000000000:address=10'd200;
		12'b001000000001:address=10'd201;
		12'b001000000010:address=10'd202;
		12'b001000000011:address=10'd203;
		12'b001000000100:address=10'd204;
		12'b001000000101:address=10'd205;
		12'b001000000110:address=10'd206;
		12'b001000000111:address=10'd207;
		12'b001000001000:address=10'd208;
		12'b001000001001:address=10'd209;
		12'b001000010000:address=10'd210;
		12'b001000010001:address=10'd211;
		12'b001000010010:address=10'd212;
		12'b001000010011:address=10'd213;
		12'b001000010100:address=10'd214;
		12'b001000010101:address=10'd215;
		12'b001000010110:address=10'd216;
		12'b001000010111:address=10'd217;
		12'b001000011000:address=10'd218;
		12'b001000011001:address=10'd219;
		12'b001000100000:address=10'd220;
		12'b001000100001:address=10'd221;
		12'b001000100010:address=10'd222;
		12'b001000100011:address=10'd223;
		12'b001000100100:address=10'd224;
		12'b001000100101:address=10'd225;
		12'b001000100110:address=10'd226;
		12'b001000100111:address=10'd227;
		12'b001000101000:address=10'd228;
		12'b001000101001:address=10'd229;
		12'b001000110000:address=10'd230;
		12'b001000110001:address=10'd231;
		12'b001000110010:address=10'd232;
		12'b001000110011:address=10'd233;
		12'b001000110100:address=10'd234;
		12'b001000110101:address=10'd235;
		12'b001000110110:address=10'd236;
		12'b001000110111:address=10'd237;
		12'b001000111000:address=10'd238;
		12'b001000111001:address=10'd239;
		12'b001001000000:address=10'd240;
		12'b001001000001:address=10'd241;
		12'b001001000010:address=10'd242;
		12'b001001000011:address=10'd243;
		12'b001001000100:address=10'd244;
		12'b001001000101:address=10'd245;
		12'b001001000110:address=10'd246;
		12'b001001000111:address=10'd247;
		12'b001001001000:address=10'd248;
		12'b001001001001:address=10'd249;
		12'b001001010000:address=10'd250;
		12'b001001010001:address=10'd251;
		12'b001001010010:address=10'd252;
		12'b001001010011:address=10'd253;
		12'b001001010100:address=10'd254;
		12'b001001010101:address=10'd255;
		12'b001001010110:address=10'd256;
		12'b001001010111:address=10'd257;
		12'b001001011000:address=10'd258;
		12'b001001011001:address=10'd259;
		12'b001001100000:address=10'd260;
		12'b001001100001:address=10'd261;
		12'b001001100010:address=10'd262;
		12'b001001100011:address=10'd263;
		12'b001001100100:address=10'd264;
		12'b001001100101:address=10'd265;
		12'b001001100110:address=10'd266;
		12'b001001100111:address=10'd267;
		12'b001001101000:address=10'd268;
		12'b001001101001:address=10'd269;
		12'b001001110000:address=10'd270;
		12'b001001110001:address=10'd271;
		12'b001001110010:address=10'd272;
		12'b001001110011:address=10'd273;
		12'b001001110100:address=10'd274;
		12'b001001110101:address=10'd275;
		12'b001001110110:address=10'd276;
		12'b001001110111:address=10'd277;
		12'b001001111000:address=10'd278;
		12'b001001111001:address=10'd279;
		12'b001010000000:address=10'd280;
		12'b001010000001:address=10'd281;
		12'b001010000010:address=10'd282;
		12'b001010000011:address=10'd283;
		12'b001010000100:address=10'd284;
		12'b001010000101:address=10'd285;
		12'b001010000110:address=10'd286;
		12'b001010000111:address=10'd287;
		12'b001010001000:address=10'd288;
		12'b001010001001:address=10'd289;
		12'b001010010000:address=10'd290;
		12'b001010010001:address=10'd291;
		12'b001010010010:address=10'd292;
		12'b001010010011:address=10'd293;
		12'b001010010100:address=10'd294;
		12'b001010010101:address=10'd295;
		12'b001010010110:address=10'd296;
		12'b001010010111:address=10'd297;
		12'b001010011000:address=10'd298;
		12'b001010011001:address=10'd299;
		12'b001100000000:address=10'd300;
		12'b001100000001:address=10'd301;
		12'b001100000010:address=10'd302;
		12'b001100000011:address=10'd303;
		12'b001100000100:address=10'd304;
		12'b001100000101:address=10'd305;
		12'b001100000110:address=10'd306;
		12'b001100000111:address=10'd307;
		12'b001100001000:address=10'd308;
		12'b001100001001:address=10'd309;
		12'b001100010000:address=10'd310;
		12'b001100010001:address=10'd311;
		12'b001100010010:address=10'd312;
		12'b001100010011:address=10'd313;
		12'b001100010100:address=10'd314;
		12'b001100010101:address=10'd315;
		12'b001100010110:address=10'd316;
		12'b001100010111:address=10'd317;
		12'b001100011000:address=10'd318;
		12'b001100011001:address=10'd319;
		12'b001100100000:address=10'd320;
		12'b001100100001:address=10'd321;
		12'b001100100010:address=10'd322;
		12'b001100100011:address=10'd323;
		12'b001100100100:address=10'd324;
		12'b001100100101:address=10'd325;
		12'b001100100110:address=10'd326;
		12'b001100100111:address=10'd327;
		12'b001100101000:address=10'd328;
		12'b001100101001:address=10'd329;
		12'b001100110000:address=10'd330;
		12'b001100110001:address=10'd331;
		12'b001100110010:address=10'd332;
		12'b001100110011:address=10'd333;
		12'b001100110100:address=10'd334;
		12'b001100110101:address=10'd335;
		12'b001100110110:address=10'd336;
		12'b001100110111:address=10'd337;
		12'b001100111000:address=10'd338;
		12'b001100111001:address=10'd339;
		12'b001101000000:address=10'd340;
		12'b001101000001:address=10'd341;
		12'b001101000010:address=10'd342;
		12'b001101000011:address=10'd343;
		12'b001101000100:address=10'd344;
		12'b001101000101:address=10'd345;
		12'b001101000110:address=10'd346;
		12'b001101000111:address=10'd347;
		12'b001101001000:address=10'd348;
		12'b001101001001:address=10'd349;
		12'b001101010000:address=10'd350;
		12'b001101010001:address=10'd351;
		12'b001101010010:address=10'd352;
		12'b001101010011:address=10'd353;
		12'b001101010100:address=10'd354;
		12'b001101010101:address=10'd355;
		12'b001101010110:address=10'd356;
		12'b001101010111:address=10'd357;
		12'b001101011000:address=10'd358;
		12'b001101011001:address=10'd359;
		12'b001101100000:address=10'd360;
		12'b001101100001:address=10'd361;
		12'b001101100010:address=10'd362;
		12'b001101100011:address=10'd363;
		12'b001101100100:address=10'd364;
		12'b001101100101:address=10'd365;
		12'b001101100110:address=10'd366;
		12'b001101100111:address=10'd367;
		12'b001101101000:address=10'd368;
		12'b001101101001:address=10'd369;
		12'b001101110000:address=10'd370;
		12'b001101110001:address=10'd371;
		12'b001101110010:address=10'd372;
		12'b001101110011:address=10'd373;
		12'b001101110100:address=10'd374;
		12'b001101110101:address=10'd375;
		12'b001101110110:address=10'd376;
		12'b001101110111:address=10'd377;
		12'b001101111000:address=10'd378;
		12'b001101111001:address=10'd379;
		12'b001110000000:address=10'd380;
		12'b001110000001:address=10'd381;
		12'b001110000010:address=10'd382;
		12'b001110000011:address=10'd383;
		12'b001110000100:address=10'd384;
		12'b001110000101:address=10'd385;
		12'b001110000110:address=10'd386;
		12'b001110000111:address=10'd387;
		12'b001110001000:address=10'd388;
		12'b001110001001:address=10'd389;
		12'b001110010000:address=10'd390;
		12'b001110010001:address=10'd391;
		12'b001110010010:address=10'd392;
		12'b001110010011:address=10'd393;
		12'b001110010100:address=10'd394;
		12'b001110010101:address=10'd395;
		12'b001110010110:address=10'd396;
		12'b001110010111:address=10'd397;
		12'b001110011000:address=10'd398;
		12'b001110011001:address=10'd399;
		12'b010000000000:address=10'd400;
		12'b010000000001:address=10'd401;
		12'b010000000010:address=10'd402;
		12'b010000000011:address=10'd403;
		12'b010000000100:address=10'd404;
		12'b010000000101:address=10'd405;
		12'b010000000110:address=10'd406;
		12'b010000000111:address=10'd407;
		12'b010000001000:address=10'd408;
		12'b010000001001:address=10'd409;
		12'b010000010000:address=10'd410;
		12'b010000010001:address=10'd411;
		12'b010000010010:address=10'd412;
		12'b010000010011:address=10'd413;
		12'b010000010100:address=10'd414;
		12'b010000010101:address=10'd415;
		12'b010000010110:address=10'd416;
		12'b010000010111:address=10'd417;
		12'b010000011000:address=10'd418;
		12'b010000011001:address=10'd419;
		12'b010000100000:address=10'd420;
		12'b010000100001:address=10'd421;
		12'b010000100010:address=10'd422;
		12'b010000100011:address=10'd423;
		12'b010000100100:address=10'd424;
		12'b010000100101:address=10'd425;
		12'b010000100110:address=10'd426;
		12'b010000100111:address=10'd427;
		12'b010000101000:address=10'd428;
		12'b010000101001:address=10'd429;
		12'b010000110000:address=10'd430;
		12'b010000110001:address=10'd431;
		12'b010000110010:address=10'd432;
		12'b010000110011:address=10'd433;
		12'b010000110100:address=10'd434;
		12'b010000110101:address=10'd435;
		12'b010000110110:address=10'd436;
		12'b010000110111:address=10'd437;
		12'b010000111000:address=10'd438;
		12'b010000111001:address=10'd439;
		12'b010001000000:address=10'd440;
		12'b010001000001:address=10'd441;
		12'b010001000010:address=10'd442;
		12'b010001000011:address=10'd443;
		12'b010001000100:address=10'd444;
		12'b010001000101:address=10'd445;
		12'b010001000110:address=10'd446;
		12'b010001000111:address=10'd447;
		12'b010001001000:address=10'd448;
		12'b010001001001:address=10'd449;
		12'b010001010000:address=10'd450;
		12'b010001010001:address=10'd451;
		12'b010001010010:address=10'd452;
		12'b010001010011:address=10'd453;
		12'b010001010100:address=10'd454;
		12'b010001010101:address=10'd455;
		12'b010001010110:address=10'd456;
		12'b010001010111:address=10'd457;
		12'b010001011000:address=10'd458;
		12'b010001011001:address=10'd459;
		12'b010001100000:address=10'd460;
		12'b010001100001:address=10'd461;
		12'b010001100010:address=10'd462;
		12'b010001100011:address=10'd463;
		12'b010001100100:address=10'd464;
		12'b010001100101:address=10'd465;
		12'b010001100110:address=10'd466;
		12'b010001100111:address=10'd467;
		12'b010001101000:address=10'd468;
		12'b010001101001:address=10'd469;
		12'b010001110000:address=10'd470;
		12'b010001110001:address=10'd471;
		12'b010001110010:address=10'd472;
		12'b010001110011:address=10'd473;
		12'b010001110100:address=10'd474;
		12'b010001110101:address=10'd475;
		12'b010001110110:address=10'd476;
		12'b010001110111:address=10'd477;
		12'b010001111000:address=10'd478;
		12'b010001111001:address=10'd479;
		12'b010010000000:address=10'd480;
		12'b010010000001:address=10'd481;
		12'b010010000010:address=10'd482;
		12'b010010000011:address=10'd483;
		12'b010010000100:address=10'd484;
		12'b010010000101:address=10'd485;
		12'b010010000110:address=10'd486;
		12'b010010000111:address=10'd487;
		12'b010010001000:address=10'd488;
		12'b010010001001:address=10'd489;
		12'b010010010000:address=10'd490;
		12'b010010010001:address=10'd491;
		12'b010010010010:address=10'd492;
		12'b010010010011:address=10'd493;
		12'b010010010100:address=10'd494;
		12'b010010010101:address=10'd495;
		12'b010010010110:address=10'd496;
		12'b010010010111:address=10'd497;
		12'b010010011000:address=10'd498;
		12'b010010011001:address=10'd499;
		12'b010100000000:address=10'd500;
		12'b010100000001:address=10'd501;
		12'b010100000010:address=10'd502;
		12'b010100000011:address=10'd503;
		12'b010100000100:address=10'd504;
		12'b010100000101:address=10'd505;
		12'b010100000110:address=10'd506;
		12'b010100000111:address=10'd507;
		12'b010100001000:address=10'd508;
		12'b010100001001:address=10'd509;
		12'b010100010000:address=10'd510;
		12'b010100010001:address=10'd511;
		12'b010100010010:address=10'd512;
		12'b010100010011:address=10'd513;
		12'b010100010100:address=10'd514;
		12'b010100010101:address=10'd515;
		12'b010100010110:address=10'd516;
		12'b010100010111:address=10'd517;
		12'b010100011000:address=10'd518;
		12'b010100011001:address=10'd519;
		12'b010100100000:address=10'd520;
		12'b010100100001:address=10'd521;
		12'b010100100010:address=10'd522;
		12'b010100100011:address=10'd523;
		12'b010100100100:address=10'd524;
		12'b010100100101:address=10'd525;
		12'b010100100110:address=10'd526;
		12'b010100100111:address=10'd527;
		12'b010100101000:address=10'd528;
		12'b010100101001:address=10'd529;
		12'b010100110000:address=10'd530;
		12'b010100110001:address=10'd531;
		12'b010100110010:address=10'd532;
		12'b010100110011:address=10'd533;
		12'b010100110100:address=10'd534;
		12'b010100110101:address=10'd535;
		12'b010100110110:address=10'd536;
		12'b010100110111:address=10'd537;
		12'b010100111000:address=10'd538;
		12'b010100111001:address=10'd539;
		12'b010101000000:address=10'd540;
		12'b010101000001:address=10'd541;
		12'b010101000010:address=10'd542;
		12'b010101000011:address=10'd543;
		12'b010101000100:address=10'd544;
		12'b010101000101:address=10'd545;
		12'b010101000110:address=10'd546;
		12'b010101000111:address=10'd547;
		12'b010101001000:address=10'd548;
		12'b010101001001:address=10'd549;
		12'b010101010000:address=10'd550;
		12'b010101010001:address=10'd551;
		12'b010101010010:address=10'd552;
		12'b010101010011:address=10'd553;
		12'b010101010100:address=10'd554;
		12'b010101010101:address=10'd555;
		12'b010101010110:address=10'd556;
		12'b010101010111:address=10'd557;
		12'b010101011000:address=10'd558;
		12'b010101011001:address=10'd559;
		12'b010101100000:address=10'd560;
		12'b010101100001:address=10'd561;
		12'b010101100010:address=10'd562;
		12'b010101100011:address=10'd563;
		12'b010101100100:address=10'd564;
		12'b010101100101:address=10'd565;
		12'b010101100110:address=10'd566;
		12'b010101100111:address=10'd567;
		12'b010101101000:address=10'd568;
		12'b010101101001:address=10'd569;
		12'b010101110000:address=10'd570;
		12'b010101110001:address=10'd571;
		12'b010101110010:address=10'd572;
		12'b010101110011:address=10'd573;
		12'b010101110100:address=10'd574;
		12'b010101110101:address=10'd575;
		12'b010101110110:address=10'd576;
		12'b010101110111:address=10'd577;
		12'b010101111000:address=10'd578;
		12'b010101111001:address=10'd579;
		12'b010110000000:address=10'd580;
		12'b010110000001:address=10'd581;
		12'b010110000010:address=10'd582;
		12'b010110000011:address=10'd583;
		12'b010110000100:address=10'd584;
		12'b010110000101:address=10'd585;
		12'b010110000110:address=10'd586;
		12'b010110000111:address=10'd587;
		12'b010110001000:address=10'd588;
		12'b010110001001:address=10'd589;
		12'b010110010000:address=10'd590;
		12'b010110010001:address=10'd591;
		12'b010110010010:address=10'd592;
		12'b010110010011:address=10'd593;
		12'b010110010100:address=10'd594;
		12'b010110010101:address=10'd595;
		12'b010110010110:address=10'd596;
		12'b010110010111:address=10'd597;
		12'b010110011000:address=10'd598;
		12'b010110011001:address=10'd599;
		12'b011000000000:address=10'd600;
		12'b011000000001:address=10'd601;
		12'b011000000010:address=10'd602;
		12'b011000000011:address=10'd603;
		12'b011000000100:address=10'd604;
		12'b011000000101:address=10'd605;
		12'b011000000110:address=10'd606;
		12'b011000000111:address=10'd607;
		12'b011000001000:address=10'd608;
		12'b011000001001:address=10'd609;
		12'b011000010000:address=10'd610;
		12'b011000010001:address=10'd611;
		12'b011000010010:address=10'd612;
		12'b011000010011:address=10'd613;
		12'b011000010100:address=10'd614;
		12'b011000010101:address=10'd615;
		12'b011000010110:address=10'd616;
		12'b011000010111:address=10'd617;
		12'b011000011000:address=10'd618;
		12'b011000011001:address=10'd619;
		12'b011000100000:address=10'd620;
		12'b011000100001:address=10'd621;
		12'b011000100010:address=10'd622;
		12'b011000100011:address=10'd623;
		12'b011000100100:address=10'd624;
		12'b011000100101:address=10'd625;
		12'b011000100110:address=10'd626;
		12'b011000100111:address=10'd627;
		12'b011000101000:address=10'd628;
		12'b011000101001:address=10'd629;
		12'b011000110000:address=10'd630;
		12'b011000110001:address=10'd631;
		12'b011000110010:address=10'd632;
		12'b011000110011:address=10'd633;
		12'b011000110100:address=10'd634;
		12'b011000110101:address=10'd635;
		12'b011000110110:address=10'd636;
		12'b011000110111:address=10'd637;
		12'b011000111000:address=10'd638;
		12'b011000111001:address=10'd639;
		12'b011001000000:address=10'd640;
		12'b011001000001:address=10'd641;
		12'b011001000010:address=10'd642;
		12'b011001000011:address=10'd643;
		12'b011001000100:address=10'd644;
		12'b011001000101:address=10'd645;
		12'b011001000110:address=10'd646;
		12'b011001000111:address=10'd647;
		12'b011001001000:address=10'd648;
		12'b011001001001:address=10'd649;
		12'b011001010000:address=10'd650;
		12'b011001010001:address=10'd651;
		12'b011001010010:address=10'd652;
		12'b011001010011:address=10'd653;
		12'b011001010100:address=10'd654;
		12'b011001010101:address=10'd655;
		12'b011001010110:address=10'd656;
		12'b011001010111:address=10'd657;
		12'b011001011000:address=10'd658;
		12'b011001011001:address=10'd659;
		12'b011001100000:address=10'd660;
		12'b011001100001:address=10'd661;
		12'b011001100010:address=10'd662;
		12'b011001100011:address=10'd663;
		12'b011001100100:address=10'd664;
		12'b011001100101:address=10'd665;
		12'b011001100110:address=10'd666;
		12'b011001100111:address=10'd667;
		12'b011001101000:address=10'd668;
		12'b011001101001:address=10'd669;
		12'b011001110000:address=10'd670;
		12'b011001110001:address=10'd671;
		12'b011001110010:address=10'd672;
		12'b011001110011:address=10'd673;
		12'b011001110100:address=10'd674;
		12'b011001110101:address=10'd675;
		12'b011001110110:address=10'd676;
		12'b011001110111:address=10'd677;
		12'b011001111000:address=10'd678;
		12'b011001111001:address=10'd679;
		12'b011010000000:address=10'd680;
		12'b011010000001:address=10'd681;
		12'b011010000010:address=10'd682;
		12'b011010000011:address=10'd683;
		12'b011010000100:address=10'd684;
		12'b011010000101:address=10'd685;
		12'b011010000110:address=10'd686;
		12'b011010000111:address=10'd687;
		12'b011010001000:address=10'd688;
		12'b011010001001:address=10'd689;
		12'b011010010000:address=10'd690;
		12'b011010010001:address=10'd691;
		12'b011010010010:address=10'd692;
		12'b011010010011:address=10'd693;
		12'b011010010100:address=10'd694;
		12'b011010010101:address=10'd695;
		12'b011010010110:address=10'd696;
		12'b011010010111:address=10'd697;
		12'b011010011000:address=10'd698;
		12'b011010011001:address=10'd699;
    endcase
end


endmodule
module testBPartCounter();
    reg trigger;
    reg SysRst;
    wire [9:0] address;
    BPartCounter U1(trigger,SysRst,address);
    initial begin
        SysRst = 1;
        trigger =1;
        #5
        SysRst =0;

    end
    always begin
        #5
        trigger = ~trigger;

    end

endmodule
