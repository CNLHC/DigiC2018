module parity(
    input [7:0]data,
    output reg paritybit
);
always@(*) begin
    case(data)
//#for i in range(0,256):
//#    bitstring = "{0:08b}".format(i)
//#    print("8'b{0:s}:parity={1:d};".format(bitstring,list(bitstring).count('1')%2))
    8'b00000000:paritybit=0;
    8'b00000001:paritybit=1;
    8'b00000010:paritybit=1;
    8'b00000011:paritybit=0;
    8'b00000100:paritybit=1;
    8'b00000101:paritybit=0;
    8'b00000110:paritybit=0;
    8'b00000111:paritybit=1;
    8'b00001000:paritybit=1;
    8'b00001001:paritybit=0;
    8'b00001010:paritybit=0;
    8'b00001011:paritybit=1;
    8'b00001100:paritybit=0;
    8'b00001101:paritybit=1;
    8'b00001110:paritybit=1;
    8'b00001111:paritybit=0;
    8'b00010000:paritybit=1;
    8'b00010001:paritybit=0;
    8'b00010010:paritybit=0;
    8'b00010011:paritybit=1;
    8'b00010100:paritybit=0;
    8'b00010101:paritybit=1;
    8'b00010110:paritybit=1;
    8'b00010111:paritybit=0;
    8'b00011000:paritybit=0;
    8'b00011001:paritybit=1;
    8'b00011010:paritybit=1;
    8'b00011011:paritybit=0;
    8'b00011100:paritybit=1;
    8'b00011101:paritybit=0;
    8'b00011110:paritybit=0;
    8'b00011111:paritybit=1;
    8'b00100000:paritybit=1;
    8'b00100001:paritybit=0;
    8'b00100010:paritybit=0;
    8'b00100011:paritybit=1;
    8'b00100100:paritybit=0;
    8'b00100101:paritybit=1;
    8'b00100110:paritybit=1;
    8'b00100111:paritybit=0;
    8'b00101000:paritybit=0;
    8'b00101001:paritybit=1;
    8'b00101010:paritybit=1;
    8'b00101011:paritybit=0;
    8'b00101100:paritybit=1;
    8'b00101101:paritybit=0;
    8'b00101110:paritybit=0;
    8'b00101111:paritybit=1;
    8'b00110000:paritybit=0;
    8'b00110001:paritybit=1;
    8'b00110010:paritybit=1;
    8'b00110011:paritybit=0;
    8'b00110100:paritybit=1;
    8'b00110101:paritybit=0;
    8'b00110110:paritybit=0;
    8'b00110111:paritybit=1;
    8'b00111000:paritybit=1;
    8'b00111001:paritybit=0;
    8'b00111010:paritybit=0;
    8'b00111011:paritybit=1;
    8'b00111100:paritybit=0;
    8'b00111101:paritybit=1;
    8'b00111110:paritybit=1;
    8'b00111111:paritybit=0;
    8'b01000000:paritybit=1;
    8'b01000001:paritybit=0;
    8'b01000010:paritybit=0;
    8'b01000011:paritybit=1;
    8'b01000100:paritybit=0;
    8'b01000101:paritybit=1;
    8'b01000110:paritybit=1;
    8'b01000111:paritybit=0;
    8'b01001000:paritybit=0;
    8'b01001001:paritybit=1;
    8'b01001010:paritybit=1;
    8'b01001011:paritybit=0;
    8'b01001100:paritybit=1;
    8'b01001101:paritybit=0;
    8'b01001110:paritybit=0;
    8'b01001111:paritybit=1;
    8'b01010000:paritybit=0;
    8'b01010001:paritybit=1;
    8'b01010010:paritybit=1;
    8'b01010011:paritybit=0;
    8'b01010100:paritybit=1;
    8'b01010101:paritybit=0;
    8'b01010110:paritybit=0;
    8'b01010111:paritybit=1;
    8'b01011000:paritybit=1;
    8'b01011001:paritybit=0;
    8'b01011010:paritybit=0;
    8'b01011011:paritybit=1;
    8'b01011100:paritybit=0;
    8'b01011101:paritybit=1;
    8'b01011110:paritybit=1;
    8'b01011111:paritybit=0;
    8'b01100000:paritybit=0;
    8'b01100001:paritybit=1;
    8'b01100010:paritybit=1;
    8'b01100011:paritybit=0;
    8'b01100100:paritybit=1;
    8'b01100101:paritybit=0;
    8'b01100110:paritybit=0;
    8'b01100111:paritybit=1;
    8'b01101000:paritybit=1;
    8'b01101001:paritybit=0;
    8'b01101010:paritybit=0;
    8'b01101011:paritybit=1;
    8'b01101100:paritybit=0;
    8'b01101101:paritybit=1;
    8'b01101110:paritybit=1;
    8'b01101111:paritybit=0;
    8'b01110000:paritybit=1;
    8'b01110001:paritybit=0;
    8'b01110010:paritybit=0;
    8'b01110011:paritybit=1;
    8'b01110100:paritybit=0;
    8'b01110101:paritybit=1;
    8'b01110110:paritybit=1;
    8'b01110111:paritybit=0;
    8'b01111000:paritybit=0;
    8'b01111001:paritybit=1;
    8'b01111010:paritybit=1;
    8'b01111011:paritybit=0;
    8'b01111100:paritybit=1;
    8'b01111101:paritybit=0;
    8'b01111110:paritybit=0;
    8'b01111111:paritybit=1;
    8'b10000000:paritybit=1;
    8'b10000001:paritybit=0;
    8'b10000010:paritybit=0;
    8'b10000011:paritybit=1;
    8'b10000100:paritybit=0;
    8'b10000101:paritybit=1;
    8'b10000110:paritybit=1;
    8'b10000111:paritybit=0;
    8'b10001000:paritybit=0;
    8'b10001001:paritybit=1;
    8'b10001010:paritybit=1;
    8'b10001011:paritybit=0;
    8'b10001100:paritybit=1;
    8'b10001101:paritybit=0;
    8'b10001110:paritybit=0;
    8'b10001111:paritybit=1;
    8'b10010000:paritybit=0;
    8'b10010001:paritybit=1;
    8'b10010010:paritybit=1;
    8'b10010011:paritybit=0;
    8'b10010100:paritybit=1;
    8'b10010101:paritybit=0;
    8'b10010110:paritybit=0;
    8'b10010111:paritybit=1;
    8'b10011000:paritybit=1;
    8'b10011001:paritybit=0;
    8'b10011010:paritybit=0;
    8'b10011011:paritybit=1;
    8'b10011100:paritybit=0;
    8'b10011101:paritybit=1;
    8'b10011110:paritybit=1;
    8'b10011111:paritybit=0;
    8'b10100000:paritybit=0;
    8'b10100001:paritybit=1;
    8'b10100010:paritybit=1;
    8'b10100011:paritybit=0;
    8'b10100100:paritybit=1;
    8'b10100101:paritybit=0;
    8'b10100110:paritybit=0;
    8'b10100111:paritybit=1;
    8'b10101000:paritybit=1;
    8'b10101001:paritybit=0;
    8'b10101010:paritybit=0;
    8'b10101011:paritybit=1;
    8'b10101100:paritybit=0;
    8'b10101101:paritybit=1;
    8'b10101110:paritybit=1;
    8'b10101111:paritybit=0;
    8'b10110000:paritybit=1;
    8'b10110001:paritybit=0;
    8'b10110010:paritybit=0;
    8'b10110011:paritybit=1;
    8'b10110100:paritybit=0;
    8'b10110101:paritybit=1;
    8'b10110110:paritybit=1;
    8'b10110111:paritybit=0;
    8'b10111000:paritybit=0;
    8'b10111001:paritybit=1;
    8'b10111010:paritybit=1;
    8'b10111011:paritybit=0;
    8'b10111100:paritybit=1;
    8'b10111101:paritybit=0;
    8'b10111110:paritybit=0;
    8'b10111111:paritybit=1;
    8'b11000000:paritybit=0;
    8'b11000001:paritybit=1;
    8'b11000010:paritybit=1;
    8'b11000011:paritybit=0;
    8'b11000100:paritybit=1;
    8'b11000101:paritybit=0;
    8'b11000110:paritybit=0;
    8'b11000111:paritybit=1;
    8'b11001000:paritybit=1;
    8'b11001001:paritybit=0;
    8'b11001010:paritybit=0;
    8'b11001011:paritybit=1;
    8'b11001100:paritybit=0;
    8'b11001101:paritybit=1;
    8'b11001110:paritybit=1;
    8'b11001111:paritybit=0;
    8'b11010000:paritybit=1;
    8'b11010001:paritybit=0;
    8'b11010010:paritybit=0;
    8'b11010011:paritybit=1;
    8'b11010100:paritybit=0;
    8'b11010101:paritybit=1;
    8'b11010110:paritybit=1;
    8'b11010111:paritybit=0;
    8'b11011000:paritybit=0;
    8'b11011001:paritybit=1;
    8'b11011010:paritybit=1;
    8'b11011011:paritybit=0;
    8'b11011100:paritybit=1;
    8'b11011101:paritybit=0;
    8'b11011110:paritybit=0;
    8'b11011111:paritybit=1;
    8'b11100000:paritybit=1;
    8'b11100001:paritybit=0;
    8'b11100010:paritybit=0;
    8'b11100011:paritybit=1;
    8'b11100100:paritybit=0;
    8'b11100101:paritybit=1;
    8'b11100110:paritybit=1;
    8'b11100111:paritybit=0;
    8'b11101000:paritybit=0;
    8'b11101001:paritybit=1;
    8'b11101010:paritybit=1;
    8'b11101011:paritybit=0;
    8'b11101100:paritybit=1;
    8'b11101101:paritybit=0;
    8'b11101110:paritybit=0;
    8'b11101111:paritybit=1;
    8'b11110000:paritybit=0;
    8'b11110001:paritybit=1;
    8'b11110010:paritybit=1;
    8'b11110011:paritybit=0;
    8'b11110100:paritybit=1;
    8'b11110101:paritybit=0;
    8'b11110110:paritybit=0;
    8'b11110111:paritybit=1;
    8'b11111000:paritybit=1;
    8'b11111001:paritybit=0;
    8'b11111010:paritybit=0;
    8'b11111011:paritybit=1;
    8'b11111100:paritybit=0;
    8'b11111101:paritybit=1;
    8'b11111110:paritybit=1;
    8'b11111111:paritybit=0;
    endcase
end
endmodule
