`timescale 1ns / 1ps
`define tubeDigit0 8'11111100
`define tubeDigit1 8'00001100
`define tubeDigit2 8'11011010
`define tubeDigit3 8'11110010
`define tubeDigit4 8'01100110
`define tubeDigit5 8'10110110
`define tubeDigit6 8'10111110
`define tubeDigit7 8'11100000
`define tubeDigit8 8'11111110
`define tubeDigit9 8'11110110
`define tubeDigitA 8'11101110
`define tubeDigitB 8'00111110
`define tubeDigitC 8'10011100
`define tubeDigitD 8'01111010
`define tubeDigitE 8'10011110
`define tubeDigitF 8'10001110
`define  DIV_COE 25000000
module tubeDriver(
	input [7:0]data,
	output [7:0]HEX);

endmodule
