module power(
    output H,
    output L);
assign H=1'b1;
assign L=1'b0;
endmodule
