module PROM1024x16(
    input  [9:0]address,
    output [15:0]word)
always @(*) begin
    case(address)begin


    endcase
end
endmodule

